// *********************************************************************
// IBM CONFIDENTIAL BACKGROUND TECHNOLOGY: VERIFICATION ENVIRONMENT FILE
// *********************************************************************

`ifndef _TL_SVH
`define _TL_SVH

`include "tl_dl_if.sv"
`include "tl_tx_driver.sv"
`include "tl_tx_monitor.sv"
`include "tl_tx_seqr.sv"
`include "tl_rx_monitor.sv"
`include "tl_agent.sv"

`endif

