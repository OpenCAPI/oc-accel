/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
`ifndef _TL_BFM_PKG_SVH_
`define _TL_BFM_PKG_SVH_

//CONFIG
//INTERFACE & TRANSACTIONS
//MANAGER
`include "../util/util.svh"

//SCOREBOARDS
`include "../sb/sb.svh"

//MONITORS
//DRIVER
//AGENTS
`include "../tl/tl.svh"

//TL BFM TOP
//`include "tl_bfm_env.sv"

//TEST LIST
`include "../seq_lib/test_list.svh"

`endif // _TL_BFM_PKG_SVH_
