/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
`define VLIB_BYPASS_POWER_CG
`define NV_FPGA_FIFOGEN
`define FPGA
`define DESIGNWARE_NOEXIST
`define NV_FPGA_SYSTEM
`define NV_FPGA_UNIT
`define XSDB_SLV_DIS
`define NV_LARGE
