// *********************************************************************
// IBM CONFIDENTIAL BACKGROUND TECHNOLOGY: VERIFICATION ENVIRONMENT FILE
// *********************************************************************

`ifndef _UTIL_SVH
`define _UTIL_SVH

`include "tl_cfg_obj.sv"
`include "tl_tx_trans.sv"
`include "tl_rx_trans.sv"
`include "dl_credit_trans.sv"
`include "host_mem_model.sv"
`include "tl_manager.sv"
`include "tl_trans.sv"

`endif

