/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
`ifndef _TEST_LIST_SVH
`define _TEST_LIST_SVH

`include "bfm_sequence_base.sv"
`include "bfm_seq_lib.sv"
`include "bfm_seq_lib_rand_resp.sv"
`include "bfm_seq_lib_rand_axi.sv"
`include "bfm_seq_lib_rand_axi_resp.sv"
`include "odma_seq_lib.sv"
`include "odma_seq_lib_unalign.sv"
`include "bfm_seq_lib_mmio_intrp.sv"

`endif
