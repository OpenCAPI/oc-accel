/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
//------------------------------------------------------------------------------
//
// CLASS: intrp_interface
//
//------------------------------------------------------------------------------
`ifndef _INTRP_INTERFACE_SV
`define _INTRP_INTERFACE_SV

interface intrp_interface (input logic action_clock, input logic action_rst_n);

    logic             intrp_req;
    logic             intrp_ack;
    logic      [63:0] intrp_src;
    logic       [8:0] intrp_ctx;

endinterface: intrp_interface

`endif
