`define NVTOOLS_SYNC2D_GENERIC_CELL
`define PRAND_OFF
