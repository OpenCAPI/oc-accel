/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
`ifndef _UTIL_SVH
`define _UTIL_SVH

`include "tl_cfg_obj.sv"
`include "tl_tx_trans.sv"
`include "tl_rx_trans.sv"
`include "dl_credit_trans.sv"
`include "host_mem_model.sv"
`include "tl_manager.sv"
`include "tl_trans.sv"

`endif

