`define SYNTHESIS
