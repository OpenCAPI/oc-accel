parameter   WRITEREG_NUMBER = 6;
parameter   [32*WRITEREG_NUMBER-1:0] PARAM_ARRAY = {32'h30,32'h28,32'h20,32'h1c,32'h14,32'h10};
