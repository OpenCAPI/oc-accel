/*
 * Copyright 2019 International Business Machines
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
`include "snap_global_vars.v"

module action_wrapper (
   input                                   ap_clk                   ,
   input                                   ap_rst_n                 ,
   output                                  interrupt                ,
   output [`INT_BITS-1:0]                  interrupt_src            ,
   output [`CTXW-1:0]                      interrupt_ctx            ,
   input                                   interrupt_ack            ,
    //
    // AXI Control Register inputterface
   input [ `AXI_LITE_AW-1 : 0]             s_axi_ctrl_reg_araddr    ,
   output                                  s_axi_ctrl_reg_arready   ,
   input                                   s_axi_ctrl_reg_arvalid   ,
   input [ `AXI_LITE_AW-1 : 0]             s_axi_ctrl_reg_awaddr    ,
   output                                  s_axi_ctrl_reg_awready   ,
   input                                   s_axi_ctrl_reg_awvalid   ,
   input                                   s_axi_ctrl_reg_bready    ,
   output [ 1 : 0]                         s_axi_ctrl_reg_bresp     ,
   output                                  s_axi_ctrl_reg_bvalid    ,
   output [ `AXI_LITE_DW-1 : 0]            s_axi_ctrl_reg_rdata     ,
   input                                   s_axi_ctrl_reg_rready    ,
   output [ 1 : 0]                         s_axi_ctrl_reg_rresp     ,
   output                                  s_axi_ctrl_reg_rvalid    ,
   input [ `AXI_LITE_DW-1 : 0]             s_axi_ctrl_reg_wdata     ,
   output                                  s_axi_ctrl_reg_wready    ,
   input [(`AXI_LITE_DW/8)-1 : 0]           s_axi_ctrl_reg_wstrb     ,
   input                                   s_axi_ctrl_reg_wvalid    ,
`ifdef ENABLE_AXI_CARD_MEM
`ifndef ENABLE_HBM
   output [ `AXI_CARD_MEM_ADDR_WIDTH-1 : 0]  m_axi_card_mem0_araddr   ,
   output [ 1 : 0]                         m_axi_card_mem0_arburst  ,
   output [ 3 : 0]                         m_axi_card_mem0_arcache  ,
   output [ `AXI_CARD_MEM_ID_WIDTH-1 : 0]    m_axi_card_mem0_arid     ,
   output [ 7 : 0]                         m_axi_card_mem0_arlen    ,
   output [ 1 : 0]                         m_axi_card_mem0_arlock   ,
   output [ 2 : 0]                         m_axi_card_mem0_arprot   ,
   output [ 3 : 0]                         m_axi_card_mem0_arqos    ,
   input                                   m_axi_card_mem0_arready  ,
   output [ 3 : 0]                         m_axi_card_mem0_arregion ,
   output [ 2 : 0]                         m_axi_card_mem0_arsize   ,
   output [ `AXI_CARD_MEM_USER_WIDTH-1 : 0] m_axi_card_mem0_aruser  ,
   output                                  m_axi_card_mem0_arvalid  ,
   output [ `AXI_CARD_MEM_ADDR_WIDTH-1 : 0]  m_axi_card_mem0_awaddr   ,
   output [ 1 : 0]                         m_axi_card_mem0_awburst  ,
   output [ 3 : 0]                         m_axi_card_mem0_awcache  ,
   output [ `AXI_CARD_MEM_ID_WIDTH-1 : 0]    m_axi_card_mem0_awid     ,
   output [ 7 : 0]                         m_axi_card_mem0_awlen    ,
   output [ 1 : 0]                         m_axi_card_mem0_awlock   ,
   output [ 2 : 0]                         m_axi_card_mem0_awprot   ,
   output [ 3 : 0]                         m_axi_card_mem0_awqos    ,
   input                                   m_axi_card_mem0_awready  ,
   output [ 3 : 0]                         m_axi_card_mem0_awregion ,
   output [ 2 : 0]                         m_axi_card_mem0_awsize   ,
   output [ `AXI_CARD_MEM_USER_WIDTH-1 : 0] m_axi_card_mem0_awuser  ,
   output                                  m_axi_card_mem0_awvalid  ,
   input [`AXI_CARD_MEM_ID_WIDTH-1 : 0]     m_axi_card_mem0_bid      ,
   output                                  m_axi_card_mem0_bready   ,
   input [ 1 : 0]                          m_axi_card_mem0_bresp    ,
   input [`AXI_CARD_MEM_USER_WIDTH-1 : 0]  m_axi_card_mem0_buser    ,
   input                                   m_axi_card_mem0_bvalid   ,
   input [`AXI_CARD_MEM_DATA_WIDTH-1 : 0]   m_axi_card_mem0_rdata    ,
   input [`AXI_CARD_MEM_ID_WIDTH-1 : 0]     m_axi_card_mem0_rid      ,
   input                                   m_axi_card_mem0_rlast    ,
   output                                  m_axi_card_mem0_rready   ,
   input [ 1 : 0]                          m_axi_card_mem0_rresp    ,
   input [ `AXI_CARD_MEM_USER_WIDTH-1 : 0] m_axi_card_mem0_ruser    ,
   input                                   m_axi_card_mem0_rvalid   ,
   output [`AXI_CARD_MEM_DATA_WIDTH-1 : 0]  m_axi_card_mem0_wdata    ,
   output                                  m_axi_card_mem0_wlast    ,
   input                                   m_axi_card_mem0_wready   ,
   output [(`AXI_CARD_MEM_DATA_WIDTH/8)-1 : 0] m_axi_card_mem0_wstrb  ,
   output [`AXI_CARD_MEM_USER_WIDTH-1 : 0] m_axi_card_mem0_wuser    ,
   output                                  m_axi_card_mem0_wvalid   ,

`else
   /* copy / paste the 45 following lines for a new interface */
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p0_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p0_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p0_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p0_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p0_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p0_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_arqos    ,
   input                                   m_axi_card_hbm_p0_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p0_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p0_aruser  ,
   output                                  m_axi_card_hbm_p0_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p0_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p0_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p0_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p0_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p0_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p0_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_awqos    ,
   input                                   m_axi_card_hbm_p0_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p0_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p0_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p0_awuser  ,
   output                                  m_axi_card_hbm_p0_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p0_bid      ,
   output                                  m_axi_card_hbm_p0_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p0_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p0_buser    ,
   input                                   m_axi_card_hbm_p0_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p0_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p0_rid      ,
   input                                   m_axi_card_hbm_p0_rlast    ,
   output                                  m_axi_card_hbm_p0_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p0_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p0_ruser    ,
   input                                   m_axi_card_hbm_p0_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p0_wdata    ,
   output                                  m_axi_card_hbm_p0_wlast    ,
   input                                   m_axi_card_hbm_p0_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p0_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p0_wuser    ,
   output                                  m_axi_card_hbm_p0_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p1_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p1_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p1_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p1_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p1_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p1_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_arqos    ,
   input                                   m_axi_card_hbm_p1_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p1_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p1_aruser  ,
   output                                  m_axi_card_hbm_p1_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p1_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p1_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p1_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p1_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p1_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p1_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_awqos    ,
   input                                   m_axi_card_hbm_p1_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p1_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p1_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p1_awuser  ,
   output                                  m_axi_card_hbm_p1_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p1_bid      ,
   output                                  m_axi_card_hbm_p1_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p1_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p1_buser    ,
   input                                   m_axi_card_hbm_p1_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p1_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p1_rid      ,
   input                                   m_axi_card_hbm_p1_rlast    ,
   output                                  m_axi_card_hbm_p1_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p1_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p1_ruser    ,
   input                                   m_axi_card_hbm_p1_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p1_wdata    ,
   output                                  m_axi_card_hbm_p1_wlast    ,
   input                                   m_axi_card_hbm_p1_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p1_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p1_wuser    ,
   output                                  m_axi_card_hbm_p1_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p2_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p2_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p2_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p2_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p2_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p2_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_arqos    ,
   input                                   m_axi_card_hbm_p2_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p2_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p2_aruser  ,
   output                                  m_axi_card_hbm_p2_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p2_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p2_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p2_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p2_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p2_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p2_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_awqos    ,
   input                                   m_axi_card_hbm_p2_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p2_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p2_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p2_awuser  ,
   output                                  m_axi_card_hbm_p2_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p2_bid      ,
   output                                  m_axi_card_hbm_p2_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p2_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p2_buser    ,
   input                                   m_axi_card_hbm_p2_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p2_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p2_rid      ,
   input                                   m_axi_card_hbm_p2_rlast    ,
   output                                  m_axi_card_hbm_p2_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p2_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p2_ruser    ,
   input                                   m_axi_card_hbm_p2_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p2_wdata    ,
   output                                  m_axi_card_hbm_p2_wlast    ,
   input                                   m_axi_card_hbm_p2_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p2_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p2_wuser    ,
   output                                  m_axi_card_hbm_p2_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p3_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p3_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p3_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p3_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p3_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p3_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_arqos    ,
   input                                   m_axi_card_hbm_p3_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p3_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p3_aruser  ,
   output                                  m_axi_card_hbm_p3_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p3_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p3_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p3_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p3_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p3_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p3_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_awqos    ,
   input                                   m_axi_card_hbm_p3_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p3_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p3_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p3_awuser  ,
   output                                  m_axi_card_hbm_p3_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p3_bid      ,
   output                                  m_axi_card_hbm_p3_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p3_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p3_buser    ,
   input                                   m_axi_card_hbm_p3_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p3_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p3_rid      ,
   input                                   m_axi_card_hbm_p3_rlast    ,
   output                                  m_axi_card_hbm_p3_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p3_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p3_ruser    ,
   input                                   m_axi_card_hbm_p3_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p3_wdata    ,
   output                                  m_axi_card_hbm_p3_wlast    ,
   input                                   m_axi_card_hbm_p3_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p3_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p3_wuser    ,
   output                                  m_axi_card_hbm_p3_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p4_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p4_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p4_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p4_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p4_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p4_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_arqos    ,
   input                                   m_axi_card_hbm_p4_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p4_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p4_aruser  ,
   output                                  m_axi_card_hbm_p4_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p4_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p4_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p4_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p4_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p4_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p4_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_awqos    ,
   input                                   m_axi_card_hbm_p4_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p4_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p4_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p4_awuser  ,
   output                                  m_axi_card_hbm_p4_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p4_bid      ,
   output                                  m_axi_card_hbm_p4_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p4_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p4_buser    ,
   input                                   m_axi_card_hbm_p4_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p4_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p4_rid      ,
   input                                   m_axi_card_hbm_p4_rlast    ,
   output                                  m_axi_card_hbm_p4_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p4_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p4_ruser    ,
   input                                   m_axi_card_hbm_p4_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p4_wdata    ,
   output                                  m_axi_card_hbm_p4_wlast    ,
   input                                   m_axi_card_hbm_p4_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p4_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p4_wuser    ,
   output                                  m_axi_card_hbm_p4_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p5_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p5_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p5_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p5_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p5_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p5_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_arqos    ,
   input                                   m_axi_card_hbm_p5_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p5_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p5_aruser  ,
   output                                  m_axi_card_hbm_p5_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p5_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p5_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p5_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p5_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p5_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p5_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_awqos    ,
   input                                   m_axi_card_hbm_p5_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p5_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p5_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p5_awuser  ,
   output                                  m_axi_card_hbm_p5_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p5_bid      ,
   output                                  m_axi_card_hbm_p5_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p5_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p5_buser    ,
   input                                   m_axi_card_hbm_p5_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p5_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p5_rid      ,
   input                                   m_axi_card_hbm_p5_rlast    ,
   output                                  m_axi_card_hbm_p5_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p5_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p5_ruser    ,
   input                                   m_axi_card_hbm_p5_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p5_wdata    ,
   output                                  m_axi_card_hbm_p5_wlast    ,
   input                                   m_axi_card_hbm_p5_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p5_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p5_wuser    ,
   output                                  m_axi_card_hbm_p5_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p6_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p6_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p6_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p6_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p6_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p6_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_arqos    ,
   input                                   m_axi_card_hbm_p6_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p6_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p6_aruser  ,
   output                                  m_axi_card_hbm_p6_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p6_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p6_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p6_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p6_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p6_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p6_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_awqos    ,
   input                                   m_axi_card_hbm_p6_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p6_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p6_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p6_awuser  ,
   output                                  m_axi_card_hbm_p6_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p6_bid      ,
   output                                  m_axi_card_hbm_p6_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p6_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p6_buser    ,
   input                                   m_axi_card_hbm_p6_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p6_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p6_rid      ,
   input                                   m_axi_card_hbm_p6_rlast    ,
   output                                  m_axi_card_hbm_p6_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p6_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p6_ruser    ,
   input                                   m_axi_card_hbm_p6_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p6_wdata    ,
   output                                  m_axi_card_hbm_p6_wlast    ,
   input                                   m_axi_card_hbm_p6_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p6_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p6_wuser    ,
   output                                  m_axi_card_hbm_p6_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p7_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p7_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p7_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p7_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p7_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p7_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_arqos    ,
   input                                   m_axi_card_hbm_p7_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p7_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p7_aruser  ,
   output                                  m_axi_card_hbm_p7_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p7_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p7_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p7_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p7_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p7_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p7_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_awqos    ,
   input                                   m_axi_card_hbm_p7_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p7_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p7_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p7_awuser  ,
   output                                  m_axi_card_hbm_p7_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p7_bid      ,
   output                                  m_axi_card_hbm_p7_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p7_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p7_buser    ,
   input                                   m_axi_card_hbm_p7_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p7_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p7_rid      ,
   input                                   m_axi_card_hbm_p7_rlast    ,
   output                                  m_axi_card_hbm_p7_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p7_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p7_ruser    ,
   input                                   m_axi_card_hbm_p7_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p7_wdata    ,
   output                                  m_axi_card_hbm_p7_wlast    ,
   input                                   m_axi_card_hbm_p7_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p7_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p7_wuser    ,
   output                                  m_axi_card_hbm_p7_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p8_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p8_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p8_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p8_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p8_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p8_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_arqos    ,
   input                                   m_axi_card_hbm_p8_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p8_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p8_aruser  ,
   output                                  m_axi_card_hbm_p8_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p8_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p8_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p8_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p8_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p8_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p8_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_awqos    ,
   input                                   m_axi_card_hbm_p8_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p8_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p8_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p8_awuser  ,
   output                                  m_axi_card_hbm_p8_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p8_bid      ,
   output                                  m_axi_card_hbm_p8_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p8_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p8_buser    ,
   input                                   m_axi_card_hbm_p8_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p8_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p8_rid      ,
   input                                   m_axi_card_hbm_p8_rlast    ,
   output                                  m_axi_card_hbm_p8_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p8_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p8_ruser    ,
   input                                   m_axi_card_hbm_p8_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p8_wdata    ,
   output                                  m_axi_card_hbm_p8_wlast    ,
   input                                   m_axi_card_hbm_p8_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p8_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p8_wuser    ,
   output                                  m_axi_card_hbm_p8_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p9_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p9_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p9_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p9_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p9_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p9_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_arqos    ,
   input                                   m_axi_card_hbm_p9_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p9_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p9_aruser  ,
   output                                  m_axi_card_hbm_p9_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p9_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p9_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p9_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p9_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p9_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p9_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_awqos    ,
   input                                   m_axi_card_hbm_p9_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p9_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p9_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p9_awuser  ,
   output                                  m_axi_card_hbm_p9_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p9_bid      ,
   output                                  m_axi_card_hbm_p9_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p9_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p9_buser    ,
   input                                   m_axi_card_hbm_p9_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p9_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p9_rid      ,
   input                                   m_axi_card_hbm_p9_rlast    ,
   output                                  m_axi_card_hbm_p9_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p9_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p9_ruser    ,
   input                                   m_axi_card_hbm_p9_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p9_wdata    ,
   output                                  m_axi_card_hbm_p9_wlast    ,
   input                                   m_axi_card_hbm_p9_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p9_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p9_wuser    ,
   output                                  m_axi_card_hbm_p9_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p10_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p10_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p10_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p10_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p10_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p10_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_arqos    ,
   input                                   m_axi_card_hbm_p10_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p10_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p10_aruser  ,
   output                                  m_axi_card_hbm_p10_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p10_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p10_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p10_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p10_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p10_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p10_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_awqos    ,
   input                                   m_axi_card_hbm_p10_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p10_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p10_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p10_awuser  ,
   output                                  m_axi_card_hbm_p10_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p10_bid      ,
   output                                  m_axi_card_hbm_p10_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p10_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p10_buser    ,
   input                                   m_axi_card_hbm_p10_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p10_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p10_rid      ,
   input                                   m_axi_card_hbm_p10_rlast    ,
   output                                  m_axi_card_hbm_p10_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p10_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p10_ruser    ,
   input                                   m_axi_card_hbm_p10_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p10_wdata    ,
   output                                  m_axi_card_hbm_p10_wlast    ,
   input                                   m_axi_card_hbm_p10_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p10_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p10_wuser    ,
   output                                  m_axi_card_hbm_p10_wvalid   ,

   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p11_araddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p11_arburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_arcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p11_arid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p11_arlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p11_arlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p11_arprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_arqos    ,
   input                                   m_axi_card_hbm_p11_arready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_arregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p11_arsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p11_aruser  ,
   output                                  m_axi_card_hbm_p11_arvalid  ,
   output [ `AXI_CARD_HBM_ADDR_WIDTH-1 : 0]  m_axi_card_hbm_p11_awaddr   ,
   output [ 1 : 0]                         m_axi_card_hbm_p11_awburst  ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_awcache  ,
   output [ `AXI_CARD_HBM_ID_WIDTH-1 : 0]    m_axi_card_hbm_p11_awid     ,
   output [ 7 : 0]                         m_axi_card_hbm_p11_awlen    ,
   output [ 1 : 0]                         m_axi_card_hbm_p11_awlock   ,
   output [ 2 : 0]                         m_axi_card_hbm_p11_awprot   ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_awqos    ,
   input                                   m_axi_card_hbm_p11_awready  ,
   output [ 3 : 0]                         m_axi_card_hbm_p11_awregion ,
   output [ 2 : 0]                         m_axi_card_hbm_p11_awsize   ,
   output [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p11_awuser  ,
   output                                  m_axi_card_hbm_p11_awvalid  ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p11_bid      ,
   output                                  m_axi_card_hbm_p11_bready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p11_bresp    ,
   input [`AXI_CARD_HBM_USER_WIDTH-1 : 0]  m_axi_card_hbm_p11_buser    ,
   input                                   m_axi_card_hbm_p11_bvalid   ,
   input [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]   m_axi_card_hbm_p11_rdata    ,
   input [`AXI_CARD_HBM_ID_WIDTH-1 : 0]     m_axi_card_hbm_p11_rid      ,
   input                                   m_axi_card_hbm_p11_rlast    ,
   output                                  m_axi_card_hbm_p11_rready   ,
   input [ 1 : 0]                          m_axi_card_hbm_p11_rresp    ,
   input [ `AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p11_ruser    ,
   input                                   m_axi_card_hbm_p11_rvalid   ,
   output [`AXI_CARD_HBM_DATA_WIDTH-1 : 0]  m_axi_card_hbm_p11_wdata    ,
   output                                  m_axi_card_hbm_p11_wlast    ,
   input                                   m_axi_card_hbm_p11_wready   ,
   output [(`AXI_CARD_HBM_DATA_WIDTH/8)-1 : 0] m_axi_card_hbm_p11_wstrb  ,
   output [`AXI_CARD_HBM_USER_WIDTH-1 : 0] m_axi_card_hbm_p11_wuser    ,
   output                                  m_axi_card_hbm_p11_wvalid   ,
`endif
`endif
    //
    // ETHERNET interface
`ifdef ENABLE_ETHERNET
`ifndef ENABLE_ETH_LOOP_BACK
// we define ethernet pins only if connected to an emac (no loopback)
   input [ 511 : 0]                        din_eth_TDATA    ,
   input                                   din_eth_TVALID   ,
   output                                  din_eth_TREADY   ,
   input [  63 : 0]                        din_eth_TKEEP    ,
   input [   0 : 0]                        din_eth_TUSER    ,
   input                                   din_eth_TLAST    ,
// Enable for ethernet TX
   output [ 511 : 0]                        dout_eth_TDATA    ,
   output                                   dout_eth_TVALID   ,
   input                                    dout_eth_TREADY   ,
   output [  63 : 0]                        dout_eth_TKEEP    ,
   output [   0 : 0]                        dout_eth_TUSER    ,
   output                                   dout_eth_TLAST    ,
   output                                   eth_reset         ,
`endif
`endif
    //
    // AXI Host Memory inputterface
   output [ `AXI_MM_AW-1 : 0]              m_axi_host_mem_araddr    ,
   output [ 1 : 0]                         m_axi_host_mem_arburst   ,
   output [ 3 : 0]                         m_axi_host_mem_arcache   ,
   output [ `IDW-1 : 0]                    m_axi_host_mem_arid      ,
   output [ 7 : 0]                         m_axi_host_mem_arlen     ,
   output [ 1 : 0]                         m_axi_host_mem_arlock    ,
   output [ 2 : 0]                         m_axi_host_mem_arprot    ,
   output [ 3 : 0]                         m_axi_host_mem_arqos     ,
   input                                   m_axi_host_mem_arready   ,
   output [ 3 : 0]                         m_axi_host_mem_arregion  ,
   output [ 2 : 0]                         m_axi_host_mem_arsize    ,
   output [ `AXI_ARUSER-1 : 0]             m_axi_host_mem_aruser    ,
   output                                  m_axi_host_mem_arvalid   ,
   output [ `AXI_MM_AW-1 : 0]              m_axi_host_mem_awaddr    ,
   output [ 1 : 0]                         m_axi_host_mem_awburst   ,
   output [ 3 : 0]                         m_axi_host_mem_awcache   ,
   output [ `IDW-1 : 0]                    m_axi_host_mem_awid      ,
   output [ 7 : 0]                         m_axi_host_mem_awlen     ,
   output [ 1 : 0]                         m_axi_host_mem_awlock    ,
   output [ 2 : 0]                         m_axi_host_mem_awprot    ,
   output [ 3 : 0]                         m_axi_host_mem_awqos     ,
   input                                   m_axi_host_mem_awready   ,
   output [ 3 : 0]                         m_axi_host_mem_awregion  ,
   output [ 2 : 0]                         m_axi_host_mem_awsize    ,
   output [`AXI_AWUSER-1 : 0]              m_axi_host_mem_awuser    ,
   output                                  m_axi_host_mem_awvalid   ,
   input [ `IDW-1 : 0]                     m_axi_host_mem_bid       ,
   output                                  m_axi_host_mem_bready    ,
   input [ 1 : 0]                          m_axi_host_mem_bresp     ,
   input [ `AXI_BUSER-1 : 0]               m_axi_host_mem_buser     ,
   input                                   m_axi_host_mem_bvalid    ,
   input [ `AXI_ACT_DW-1 : 0]              m_axi_host_mem_rdata     ,
   input [ `IDW-1 : 0]                     m_axi_host_mem_rid       ,
   input                                   m_axi_host_mem_rlast     ,
   output                                  m_axi_host_mem_rready    ,
   input [ 1 : 0]                          m_axi_host_mem_rresp     ,
   input [ `AXI_RUSER-1 : 0]               m_axi_host_mem_ruser     ,
   input                                   m_axi_host_mem_rvalid    ,
   output [ `AXI_ACT_DW-1 : 0]             m_axi_host_mem_wdata     ,
   output                                  m_axi_host_mem_wlast     ,
   input                                   m_axi_host_mem_wready    ,
   output [(`AXI_ACT_DW/8)-1 : 0]          m_axi_host_mem_wstrb     ,
   output [ `AXI_WUSER-1 : 0]              m_axi_host_mem_wuser     ,
   output                                  m_axi_host_mem_wvalid
    );


parameter ADDR_ACTION_TYPE = 32'h10;
parameter ADDR_RELEASE_LEVEL = 32'h14;
parameter ADDR_ACTION_INTERRUPT_SRC_ADDR_LO = 32'h18;
parameter ADDR_ACTION_INTERRUPT_SRC_ADDR_HI = 32'h1C;

reg context_q;
reg [31:0] interrupt_src_hi;
reg [31:0] interrupt_src_lo;
reg interrupt_q;
reg interrupt_wait_ack_q;
reg hls_rst_n_q;
wire interrupt_i;
wire [63:0] temp_card_mem0_araddr;
wire [63:0] temp_card_mem0_awaddr;
wire [63:0] temp_card_hbm_p0_araddr;
wire [63:0] temp_card_hbm_p0_awaddr;
wire [63:0] temp_card_hbm_p1_araddr;
wire [63:0] temp_card_hbm_p1_awaddr;
wire [63:0] temp_card_hbm_p2_araddr;
wire [63:0] temp_card_hbm_p2_awaddr;
wire [63:0] temp_card_hbm_p3_araddr;
wire [63:0] temp_card_hbm_p3_awaddr;
wire [63:0] temp_card_hbm_p4_araddr;
wire [63:0] temp_card_hbm_p4_awaddr;
wire [63:0] temp_card_hbm_p5_araddr;
wire [63:0] temp_card_hbm_p5_awaddr;
wire [63:0] temp_card_hbm_p6_araddr;
wire [63:0] temp_card_hbm_p6_awaddr;
wire [63:0] temp_card_hbm_p7_araddr;
wire [63:0] temp_card_hbm_p7_awaddr;
wire [63:0] temp_card_hbm_p8_araddr;
wire [63:0] temp_card_hbm_p8_awaddr;
wire [63:0] temp_card_hbm_p9_araddr;
wire [63:0] temp_card_hbm_p9_awaddr;
wire [63:0] temp_card_hbm_p10_araddr;
wire [63:0] temp_card_hbm_p10_awaddr;
wire [63:0] temp_card_hbm_p11_araddr;
wire [63:0] temp_card_hbm_p11_awaddr;

    // ETHERNET interface
    // we define the ethernet wrap signals only if ethernet loop back
`ifdef ENABLE_ETHERNET
`ifdef ENABLE_ETH_LOOP_BACK
wire [511:0] dwrap_eth_TDATA;
wire dwrap_eth_TVALID;
wire dwrap_eth_TREADY;
wire [63:0] dwrap_eth_TKEEP;
wire [0:0] dwrap_eth_TUSER;
wire [0:0] dwrap_eth_TLAST;
`endif
`endif



reg  [31:0] reg_rdata_hijack; //This will be ORed with the return data of hls_action
wire [31:0] temp_s_axi_ctrl_reg_rdata;

 hls_action hls_action_0 (
    .ap_clk                       ( ap_clk                  ) ,
    .ap_rst_n                     ( hls_rst_n_q             ) ,
`ifdef ENABLE_AXI_CARD_MEM
`ifndef ENABLE_HBM
    .m_axi_card_mem0_araddr       (temp_card_mem0_araddr    ) ,
    .m_axi_card_mem0_arburst      (m_axi_card_mem0_arburst  ) ,
    .m_axi_card_mem0_arcache      (m_axi_card_mem0_arcache  ) ,
    .m_axi_card_mem0_arid         (m_axi_card_mem0_arid[0]  ) ,//SR# 10394170
    .m_axi_card_mem0_arlen        (m_axi_card_mem0_arlen    ) ,
    .m_axi_card_mem0_arlock       (m_axi_card_mem0_arlock   ) ,
    .m_axi_card_mem0_arprot       (m_axi_card_mem0_arprot   ) ,
    .m_axi_card_mem0_arqos        (m_axi_card_mem0_arqos    ) ,
    .m_axi_card_mem0_arready      (m_axi_card_mem0_arready  ) ,
    .m_axi_card_mem0_arregion     (m_axi_card_mem0_arregion ) ,
    .m_axi_card_mem0_arsize       (m_axi_card_mem0_arsize   ) ,
    .m_axi_card_mem0_aruser       (m_axi_card_mem0_aruser   ) ,
    .m_axi_card_mem0_arvalid      (m_axi_card_mem0_arvalid  ) ,
    .m_axi_card_mem0_awaddr       (temp_card_mem0_awaddr    ) ,
    .m_axi_card_mem0_awburst      (m_axi_card_mem0_awburst  ) ,
    .m_axi_card_mem0_awcache      (m_axi_card_mem0_awcache  ) ,
    .m_axi_card_mem0_awid         (m_axi_card_mem0_awid[0]  ) ,//SR# 10394170
    .m_axi_card_mem0_awlen        (m_axi_card_mem0_awlen    ) ,
    .m_axi_card_mem0_awlock       (m_axi_card_mem0_awlock   ) ,
    .m_axi_card_mem0_awprot       (m_axi_card_mem0_awprot   ) ,
    .m_axi_card_mem0_awqos        (m_axi_card_mem0_awqos    ) ,
    .m_axi_card_mem0_awready      (m_axi_card_mem0_awready  ) ,
    .m_axi_card_mem0_awregion     (m_axi_card_mem0_awregion ) ,
    .m_axi_card_mem0_awsize       (m_axi_card_mem0_awsize   ) ,
    .m_axi_card_mem0_awuser       (m_axi_card_mem0_awuser   ) ,
    .m_axi_card_mem0_awvalid      (m_axi_card_mem0_awvalid  ) ,
    .m_axi_card_mem0_bid          (m_axi_card_mem0_bid[0]   ) ,//SR# 10394170
    .m_axi_card_mem0_bready       (m_axi_card_mem0_bready   ) ,
    .m_axi_card_mem0_bresp        (m_axi_card_mem0_bresp    ) ,
    .m_axi_card_mem0_buser        (m_axi_card_mem0_buser    ) ,
    .m_axi_card_mem0_bvalid       (m_axi_card_mem0_bvalid   ) ,
    .m_axi_card_mem0_rdata        (m_axi_card_mem0_rdata    ) ,
    .m_axi_card_mem0_rid          (m_axi_card_mem0_rid[0]   ) ,//SR# 10394170
    .m_axi_card_mem0_rlast        (m_axi_card_mem0_rlast    ) ,
    .m_axi_card_mem0_rready       (m_axi_card_mem0_rready   ) ,
    .m_axi_card_mem0_rresp        (m_axi_card_mem0_rresp    ) ,
    .m_axi_card_mem0_ruser        (m_axi_card_mem0_ruser    ) ,
    .m_axi_card_mem0_rvalid       (m_axi_card_mem0_rvalid   ) ,
    .m_axi_card_mem0_wdata        (m_axi_card_mem0_wdata    ) ,
    .m_axi_card_mem0_wid          (                         ) ,
    .m_axi_card_mem0_wlast        (m_axi_card_mem0_wlast    ) ,
    .m_axi_card_mem0_wready       (m_axi_card_mem0_wready   ) ,
    .m_axi_card_mem0_wstrb        (m_axi_card_mem0_wstrb    ) ,
    .m_axi_card_mem0_wuser        (m_axi_card_mem0_wuser    ) ,
    .m_axi_card_mem0_wvalid       (m_axi_card_mem0_wvalid   ) ,
`else
    /* copy / paste the 46 folloing lines to have a new HBM interface */
    .m_axi_card_hbm_p0_araddr       (temp_card_hbm_p0_araddr    ) ,
    .m_axi_card_hbm_p0_arburst      (m_axi_card_hbm_p0_arburst  ) ,
    .m_axi_card_hbm_p0_arcache      (m_axi_card_hbm_p0_arcache  ) ,
    .m_axi_card_hbm_p0_arid         (m_axi_card_hbm_p0_arid     ) ,
    .m_axi_card_hbm_p0_arlen        (m_axi_card_hbm_p0_arlen    ) ,
    .m_axi_card_hbm_p0_arlock       (m_axi_card_hbm_p0_arlock   ) ,
    .m_axi_card_hbm_p0_arprot       (m_axi_card_hbm_p0_arprot   ) ,
    .m_axi_card_hbm_p0_arqos        (m_axi_card_hbm_p0_arqos    ) ,
    .m_axi_card_hbm_p0_arready      (m_axi_card_hbm_p0_arready  ) ,
    .m_axi_card_hbm_p0_arregion     (m_axi_card_hbm_p0_arregion ) ,
    .m_axi_card_hbm_p0_arsize       (m_axi_card_hbm_p0_arsize   ) ,
    .m_axi_card_hbm_p0_aruser       (m_axi_card_hbm_p0_aruser   ) ,
    .m_axi_card_hbm_p0_arvalid      (m_axi_card_hbm_p0_arvalid  ) ,
    .m_axi_card_hbm_p0_awaddr       (temp_card_hbm_p0_awaddr    ) ,
    .m_axi_card_hbm_p0_awburst      (m_axi_card_hbm_p0_awburst  ) ,
    .m_axi_card_hbm_p0_awcache      (m_axi_card_hbm_p0_awcache  ) ,
    .m_axi_card_hbm_p0_awid         (m_axi_card_hbm_p0_awid     ) ,
    .m_axi_card_hbm_p0_awlen        (m_axi_card_hbm_p0_awlen    ) ,
    .m_axi_card_hbm_p0_awlock       (m_axi_card_hbm_p0_awlock   ) ,
    .m_axi_card_hbm_p0_awprot       (m_axi_card_hbm_p0_awprot   ) ,
    .m_axi_card_hbm_p0_awqos        (m_axi_card_hbm_p0_awqos    ) ,
    .m_axi_card_hbm_p0_awready      (m_axi_card_hbm_p0_awready  ) ,
    .m_axi_card_hbm_p0_awregion     (m_axi_card_hbm_p0_awregion ) ,
    .m_axi_card_hbm_p0_awsize       (m_axi_card_hbm_p0_awsize   ) ,
    .m_axi_card_hbm_p0_awuser       (m_axi_card_hbm_p0_awuser   ) ,
    .m_axi_card_hbm_p0_awvalid      (m_axi_card_hbm_p0_awvalid  ) ,
    .m_axi_card_hbm_p0_bid          (m_axi_card_hbm_p0_bid      ) ,
    .m_axi_card_hbm_p0_bready       (m_axi_card_hbm_p0_bready   ) ,
    .m_axi_card_hbm_p0_bresp        (m_axi_card_hbm_p0_bresp    ) ,
    .m_axi_card_hbm_p0_buser        (m_axi_card_hbm_p0_buser    ) ,
    .m_axi_card_hbm_p0_bvalid       (m_axi_card_hbm_p0_bvalid   ) ,
    .m_axi_card_hbm_p0_rdata        (m_axi_card_hbm_p0_rdata    ) ,
    .m_axi_card_hbm_p0_rid          (m_axi_card_hbm_p0_rid      ) ,
    .m_axi_card_hbm_p0_rlast        (m_axi_card_hbm_p0_rlast    ) ,
    .m_axi_card_hbm_p0_rready       (m_axi_card_hbm_p0_rready   ) ,
    .m_axi_card_hbm_p0_rresp        (m_axi_card_hbm_p0_rresp    ) ,
    .m_axi_card_hbm_p0_ruser        (m_axi_card_hbm_p0_ruser    ) ,
    .m_axi_card_hbm_p0_rvalid       (m_axi_card_hbm_p0_rvalid   ) ,
    .m_axi_card_hbm_p0_wdata        (m_axi_card_hbm_p0_wdata    ) ,
    .m_axi_card_hbm_p0_wid          (                           ) ,
    .m_axi_card_hbm_p0_wlast        (m_axi_card_hbm_p0_wlast    ) ,
    .m_axi_card_hbm_p0_wready       (m_axi_card_hbm_p0_wready   ) ,
    .m_axi_card_hbm_p0_wstrb        (m_axi_card_hbm_p0_wstrb    ) ,
    .m_axi_card_hbm_p0_wuser        (m_axi_card_hbm_p0_wuser    ) ,
    .m_axi_card_hbm_p0_wvalid       (m_axi_card_hbm_p0_wvalid   ) ,

    .m_axi_card_hbm_p1_araddr       (temp_card_hbm_p1_araddr    ) ,
    .m_axi_card_hbm_p1_arburst      (m_axi_card_hbm_p1_arburst  ) ,
    .m_axi_card_hbm_p1_arcache      (m_axi_card_hbm_p1_arcache  ) ,
    .m_axi_card_hbm_p1_arid         (m_axi_card_hbm_p1_arid     ) ,
    .m_axi_card_hbm_p1_arlen        (m_axi_card_hbm_p1_arlen    ) ,
    .m_axi_card_hbm_p1_arlock       (m_axi_card_hbm_p1_arlock   ) ,
    .m_axi_card_hbm_p1_arprot       (m_axi_card_hbm_p1_arprot   ) ,
    .m_axi_card_hbm_p1_arqos        (m_axi_card_hbm_p1_arqos    ) ,
    .m_axi_card_hbm_p1_arready      (m_axi_card_hbm_p1_arready  ) ,
    .m_axi_card_hbm_p1_arregion     (m_axi_card_hbm_p1_arregion ) ,
    .m_axi_card_hbm_p1_arsize       (m_axi_card_hbm_p1_arsize   ) ,
    .m_axi_card_hbm_p1_aruser       (m_axi_card_hbm_p1_aruser   ) ,
    .m_axi_card_hbm_p1_arvalid      (m_axi_card_hbm_p1_arvalid  ) ,
    .m_axi_card_hbm_p1_awaddr       (temp_card_hbm_p1_awaddr    ) ,
    .m_axi_card_hbm_p1_awburst      (m_axi_card_hbm_p1_awburst  ) ,
    .m_axi_card_hbm_p1_awcache      (m_axi_card_hbm_p1_awcache  ) ,
    .m_axi_card_hbm_p1_awid         (m_axi_card_hbm_p1_awid     ) ,
    .m_axi_card_hbm_p1_awlen        (m_axi_card_hbm_p1_awlen    ) ,
    .m_axi_card_hbm_p1_awlock       (m_axi_card_hbm_p1_awlock   ) ,
    .m_axi_card_hbm_p1_awprot       (m_axi_card_hbm_p1_awprot   ) ,
    .m_axi_card_hbm_p1_awqos        (m_axi_card_hbm_p1_awqos    ) ,
    .m_axi_card_hbm_p1_awready      (m_axi_card_hbm_p1_awready  ) ,
    .m_axi_card_hbm_p1_awregion     (m_axi_card_hbm_p1_awregion ) ,
    .m_axi_card_hbm_p1_awsize       (m_axi_card_hbm_p1_awsize   ) ,
    .m_axi_card_hbm_p1_awuser       (m_axi_card_hbm_p1_awuser   ) ,
    .m_axi_card_hbm_p1_awvalid      (m_axi_card_hbm_p1_awvalid  ) ,
    .m_axi_card_hbm_p1_bid          (m_axi_card_hbm_p1_bid      ) ,
    .m_axi_card_hbm_p1_bready       (m_axi_card_hbm_p1_bready   ) ,
    .m_axi_card_hbm_p1_bresp        (m_axi_card_hbm_p1_bresp    ) ,
    .m_axi_card_hbm_p1_buser        (m_axi_card_hbm_p1_buser    ) ,
    .m_axi_card_hbm_p1_bvalid       (m_axi_card_hbm_p1_bvalid   ) ,
    .m_axi_card_hbm_p1_rdata        (m_axi_card_hbm_p1_rdata    ) ,
    .m_axi_card_hbm_p1_rid          (m_axi_card_hbm_p1_rid      ) ,
    .m_axi_card_hbm_p1_rlast        (m_axi_card_hbm_p1_rlast    ) ,
    .m_axi_card_hbm_p1_rready       (m_axi_card_hbm_p1_rready   ) ,
    .m_axi_card_hbm_p1_rresp        (m_axi_card_hbm_p1_rresp    ) ,
    .m_axi_card_hbm_p1_ruser        (m_axi_card_hbm_p1_ruser    ) ,
    .m_axi_card_hbm_p1_rvalid       (m_axi_card_hbm_p1_rvalid   ) ,
    .m_axi_card_hbm_p1_wdata        (m_axi_card_hbm_p1_wdata    ) ,
    .m_axi_card_hbm_p1_wid          (                           ) ,
    .m_axi_card_hbm_p1_wlast        (m_axi_card_hbm_p1_wlast    ) ,
    .m_axi_card_hbm_p1_wready       (m_axi_card_hbm_p1_wready   ) ,
    .m_axi_card_hbm_p1_wstrb        (m_axi_card_hbm_p1_wstrb    ) ,
    .m_axi_card_hbm_p1_wuser        (m_axi_card_hbm_p1_wuser    ) ,
    .m_axi_card_hbm_p1_wvalid       (m_axi_card_hbm_p1_wvalid   ) ,

    .m_axi_card_hbm_p2_araddr       (temp_card_hbm_p2_araddr    ) ,
    .m_axi_card_hbm_p2_arburst      (m_axi_card_hbm_p2_arburst  ) ,
    .m_axi_card_hbm_p2_arcache      (m_axi_card_hbm_p2_arcache  ) ,
    .m_axi_card_hbm_p2_arid         (m_axi_card_hbm_p2_arid     ) ,
    .m_axi_card_hbm_p2_arlen        (m_axi_card_hbm_p2_arlen    ) ,
    .m_axi_card_hbm_p2_arlock       (m_axi_card_hbm_p2_arlock   ) ,
    .m_axi_card_hbm_p2_arprot       (m_axi_card_hbm_p2_arprot   ) ,
    .m_axi_card_hbm_p2_arqos        (m_axi_card_hbm_p2_arqos    ) ,
    .m_axi_card_hbm_p2_arready      (m_axi_card_hbm_p2_arready  ) ,
    .m_axi_card_hbm_p2_arregion     (m_axi_card_hbm_p2_arregion ) ,
    .m_axi_card_hbm_p2_arsize       (m_axi_card_hbm_p2_arsize   ) ,
    .m_axi_card_hbm_p2_aruser       (m_axi_card_hbm_p2_aruser   ) ,
    .m_axi_card_hbm_p2_arvalid      (m_axi_card_hbm_p2_arvalid  ) ,
    .m_axi_card_hbm_p2_awaddr       (temp_card_hbm_p2_awaddr    ) ,
    .m_axi_card_hbm_p2_awburst      (m_axi_card_hbm_p2_awburst  ) ,
    .m_axi_card_hbm_p2_awcache      (m_axi_card_hbm_p2_awcache  ) ,
    .m_axi_card_hbm_p2_awid         (m_axi_card_hbm_p2_awid     ) ,
    .m_axi_card_hbm_p2_awlen        (m_axi_card_hbm_p2_awlen    ) ,
    .m_axi_card_hbm_p2_awlock       (m_axi_card_hbm_p2_awlock   ) ,
    .m_axi_card_hbm_p2_awprot       (m_axi_card_hbm_p2_awprot   ) ,
    .m_axi_card_hbm_p2_awqos        (m_axi_card_hbm_p2_awqos    ) ,
    .m_axi_card_hbm_p2_awready      (m_axi_card_hbm_p2_awready  ) ,
    .m_axi_card_hbm_p2_awregion     (m_axi_card_hbm_p2_awregion ) ,
    .m_axi_card_hbm_p2_awsize       (m_axi_card_hbm_p2_awsize   ) ,
    .m_axi_card_hbm_p2_awuser       (m_axi_card_hbm_p2_awuser   ) ,
    .m_axi_card_hbm_p2_awvalid      (m_axi_card_hbm_p2_awvalid  ) ,
    .m_axi_card_hbm_p2_bid          (m_axi_card_hbm_p2_bid      ) ,
    .m_axi_card_hbm_p2_bready       (m_axi_card_hbm_p2_bready   ) ,
    .m_axi_card_hbm_p2_bresp        (m_axi_card_hbm_p2_bresp    ) ,
    .m_axi_card_hbm_p2_buser        (m_axi_card_hbm_p2_buser    ) ,
    .m_axi_card_hbm_p2_bvalid       (m_axi_card_hbm_p2_bvalid   ) ,
    .m_axi_card_hbm_p2_rdata        (m_axi_card_hbm_p2_rdata    ) ,
    .m_axi_card_hbm_p2_rid          (m_axi_card_hbm_p2_rid      ) ,
    .m_axi_card_hbm_p2_rlast        (m_axi_card_hbm_p2_rlast    ) ,
    .m_axi_card_hbm_p2_rready       (m_axi_card_hbm_p2_rready   ) ,
    .m_axi_card_hbm_p2_rresp        (m_axi_card_hbm_p2_rresp    ) ,
    .m_axi_card_hbm_p2_ruser        (m_axi_card_hbm_p2_ruser    ) ,
    .m_axi_card_hbm_p2_rvalid       (m_axi_card_hbm_p2_rvalid   ) ,
    .m_axi_card_hbm_p2_wdata        (m_axi_card_hbm_p2_wdata    ) ,
    .m_axi_card_hbm_p2_wid          (                           ) ,
    .m_axi_card_hbm_p2_wlast        (m_axi_card_hbm_p2_wlast    ) ,
    .m_axi_card_hbm_p2_wready       (m_axi_card_hbm_p2_wready   ) ,
    .m_axi_card_hbm_p2_wstrb        (m_axi_card_hbm_p2_wstrb    ) ,
    .m_axi_card_hbm_p2_wuser        (m_axi_card_hbm_p2_wuser    ) ,
    .m_axi_card_hbm_p2_wvalid       (m_axi_card_hbm_p2_wvalid   ) ,

    .m_axi_card_hbm_p3_araddr       (temp_card_hbm_p3_araddr    ) ,
    .m_axi_card_hbm_p3_arburst      (m_axi_card_hbm_p3_arburst  ) ,
    .m_axi_card_hbm_p3_arcache      (m_axi_card_hbm_p3_arcache  ) ,
    .m_axi_card_hbm_p3_arid         (m_axi_card_hbm_p3_arid     ) ,
    .m_axi_card_hbm_p3_arlen        (m_axi_card_hbm_p3_arlen    ) ,
    .m_axi_card_hbm_p3_arlock       (m_axi_card_hbm_p3_arlock   ) ,
    .m_axi_card_hbm_p3_arprot       (m_axi_card_hbm_p3_arprot   ) ,
    .m_axi_card_hbm_p3_arqos        (m_axi_card_hbm_p3_arqos    ) ,
    .m_axi_card_hbm_p3_arready      (m_axi_card_hbm_p3_arready  ) ,
    .m_axi_card_hbm_p3_arregion     (m_axi_card_hbm_p3_arregion ) ,
    .m_axi_card_hbm_p3_arsize       (m_axi_card_hbm_p3_arsize   ) ,
    .m_axi_card_hbm_p3_aruser       (m_axi_card_hbm_p3_aruser   ) ,
    .m_axi_card_hbm_p3_arvalid      (m_axi_card_hbm_p3_arvalid  ) ,
    .m_axi_card_hbm_p3_awaddr       (temp_card_hbm_p3_awaddr    ) ,
    .m_axi_card_hbm_p3_awburst      (m_axi_card_hbm_p3_awburst  ) ,
    .m_axi_card_hbm_p3_awcache      (m_axi_card_hbm_p3_awcache  ) ,
    .m_axi_card_hbm_p3_awid         (m_axi_card_hbm_p3_awid     ) ,
    .m_axi_card_hbm_p3_awlen        (m_axi_card_hbm_p3_awlen    ) ,
    .m_axi_card_hbm_p3_awlock       (m_axi_card_hbm_p3_awlock   ) ,
    .m_axi_card_hbm_p3_awprot       (m_axi_card_hbm_p3_awprot   ) ,
    .m_axi_card_hbm_p3_awqos        (m_axi_card_hbm_p3_awqos    ) ,
    .m_axi_card_hbm_p3_awready      (m_axi_card_hbm_p3_awready  ) ,
    .m_axi_card_hbm_p3_awregion     (m_axi_card_hbm_p3_awregion ) ,
    .m_axi_card_hbm_p3_awsize       (m_axi_card_hbm_p3_awsize   ) ,
    .m_axi_card_hbm_p3_awuser       (m_axi_card_hbm_p3_awuser   ) ,
    .m_axi_card_hbm_p3_awvalid      (m_axi_card_hbm_p3_awvalid  ) ,
    .m_axi_card_hbm_p3_bid          (m_axi_card_hbm_p3_bid      ) ,
    .m_axi_card_hbm_p3_bready       (m_axi_card_hbm_p3_bready   ) ,
    .m_axi_card_hbm_p3_bresp        (m_axi_card_hbm_p3_bresp    ) ,
    .m_axi_card_hbm_p3_buser        (m_axi_card_hbm_p3_buser    ) ,
    .m_axi_card_hbm_p3_bvalid       (m_axi_card_hbm_p3_bvalid   ) ,
    .m_axi_card_hbm_p3_rdata        (m_axi_card_hbm_p3_rdata    ) ,
    .m_axi_card_hbm_p3_rid          (m_axi_card_hbm_p3_rid      ) ,
    .m_axi_card_hbm_p3_rlast        (m_axi_card_hbm_p3_rlast    ) ,
    .m_axi_card_hbm_p3_rready       (m_axi_card_hbm_p3_rready   ) ,
    .m_axi_card_hbm_p3_rresp        (m_axi_card_hbm_p3_rresp    ) ,
    .m_axi_card_hbm_p3_ruser        (m_axi_card_hbm_p3_ruser    ) ,
    .m_axi_card_hbm_p3_rvalid       (m_axi_card_hbm_p3_rvalid   ) ,
    .m_axi_card_hbm_p3_wdata        (m_axi_card_hbm_p3_wdata    ) ,
    .m_axi_card_hbm_p3_wid          (                           ) ,
    .m_axi_card_hbm_p3_wlast        (m_axi_card_hbm_p3_wlast    ) ,
    .m_axi_card_hbm_p3_wready       (m_axi_card_hbm_p3_wready   ) ,
    .m_axi_card_hbm_p3_wstrb        (m_axi_card_hbm_p3_wstrb    ) ,
    .m_axi_card_hbm_p3_wuser        (m_axi_card_hbm_p3_wuser    ) ,
    .m_axi_card_hbm_p3_wvalid       (m_axi_card_hbm_p3_wvalid   ) ,

    .m_axi_card_hbm_p4_araddr       (temp_card_hbm_p4_araddr    ) ,
    .m_axi_card_hbm_p4_arburst      (m_axi_card_hbm_p4_arburst  ) ,
    .m_axi_card_hbm_p4_arcache      (m_axi_card_hbm_p4_arcache  ) ,
    .m_axi_card_hbm_p4_arid         (m_axi_card_hbm_p4_arid     ) ,
    .m_axi_card_hbm_p4_arlen        (m_axi_card_hbm_p4_arlen    ) ,
    .m_axi_card_hbm_p4_arlock       (m_axi_card_hbm_p4_arlock   ) ,
    .m_axi_card_hbm_p4_arprot       (m_axi_card_hbm_p4_arprot   ) ,
    .m_axi_card_hbm_p4_arqos        (m_axi_card_hbm_p4_arqos    ) ,
    .m_axi_card_hbm_p4_arready      (m_axi_card_hbm_p4_arready  ) ,
    .m_axi_card_hbm_p4_arregion     (m_axi_card_hbm_p4_arregion ) ,
    .m_axi_card_hbm_p4_arsize       (m_axi_card_hbm_p4_arsize   ) ,
    .m_axi_card_hbm_p4_aruser       (m_axi_card_hbm_p4_aruser   ) ,
    .m_axi_card_hbm_p4_arvalid      (m_axi_card_hbm_p4_arvalid  ) ,
    .m_axi_card_hbm_p4_awaddr       (temp_card_hbm_p4_awaddr    ) ,
    .m_axi_card_hbm_p4_awburst      (m_axi_card_hbm_p4_awburst  ) ,
    .m_axi_card_hbm_p4_awcache      (m_axi_card_hbm_p4_awcache  ) ,
    .m_axi_card_hbm_p4_awid         (m_axi_card_hbm_p4_awid     ) ,
    .m_axi_card_hbm_p4_awlen        (m_axi_card_hbm_p4_awlen    ) ,
    .m_axi_card_hbm_p4_awlock       (m_axi_card_hbm_p4_awlock   ) ,
    .m_axi_card_hbm_p4_awprot       (m_axi_card_hbm_p4_awprot   ) ,
    .m_axi_card_hbm_p4_awqos        (m_axi_card_hbm_p4_awqos    ) ,
    .m_axi_card_hbm_p4_awready      (m_axi_card_hbm_p4_awready  ) ,
    .m_axi_card_hbm_p4_awregion     (m_axi_card_hbm_p4_awregion ) ,
    .m_axi_card_hbm_p4_awsize       (m_axi_card_hbm_p4_awsize   ) ,
    .m_axi_card_hbm_p4_awuser       (m_axi_card_hbm_p4_awuser   ) ,
    .m_axi_card_hbm_p4_awvalid      (m_axi_card_hbm_p4_awvalid  ) ,
    .m_axi_card_hbm_p4_bid          (m_axi_card_hbm_p4_bid      ) ,
    .m_axi_card_hbm_p4_bready       (m_axi_card_hbm_p4_bready   ) ,
    .m_axi_card_hbm_p4_bresp        (m_axi_card_hbm_p4_bresp    ) ,
    .m_axi_card_hbm_p4_buser        (m_axi_card_hbm_p4_buser    ) ,
    .m_axi_card_hbm_p4_bvalid       (m_axi_card_hbm_p4_bvalid   ) ,
    .m_axi_card_hbm_p4_rdata        (m_axi_card_hbm_p4_rdata    ) ,
    .m_axi_card_hbm_p4_rid          (m_axi_card_hbm_p4_rid      ) ,
    .m_axi_card_hbm_p4_rlast        (m_axi_card_hbm_p4_rlast    ) ,
    .m_axi_card_hbm_p4_rready       (m_axi_card_hbm_p4_rready   ) ,
    .m_axi_card_hbm_p4_rresp        (m_axi_card_hbm_p4_rresp    ) ,
    .m_axi_card_hbm_p4_ruser        (m_axi_card_hbm_p4_ruser    ) ,
    .m_axi_card_hbm_p4_rvalid       (m_axi_card_hbm_p4_rvalid   ) ,
    .m_axi_card_hbm_p4_wdata        (m_axi_card_hbm_p4_wdata    ) ,
    .m_axi_card_hbm_p4_wid          (                           ) ,
    .m_axi_card_hbm_p4_wlast        (m_axi_card_hbm_p4_wlast    ) ,
    .m_axi_card_hbm_p4_wready       (m_axi_card_hbm_p4_wready   ) ,
    .m_axi_card_hbm_p4_wstrb        (m_axi_card_hbm_p4_wstrb    ) ,
    .m_axi_card_hbm_p4_wuser        (m_axi_card_hbm_p4_wuser    ) ,
    .m_axi_card_hbm_p4_wvalid       (m_axi_card_hbm_p4_wvalid   ) ,

    .m_axi_card_hbm_p5_araddr       (temp_card_hbm_p5_araddr    ) ,
    .m_axi_card_hbm_p5_arburst      (m_axi_card_hbm_p5_arburst  ) ,
    .m_axi_card_hbm_p5_arcache      (m_axi_card_hbm_p5_arcache  ) ,
    .m_axi_card_hbm_p5_arid         (m_axi_card_hbm_p5_arid     ) ,
    .m_axi_card_hbm_p5_arlen        (m_axi_card_hbm_p5_arlen    ) ,
    .m_axi_card_hbm_p5_arlock       (m_axi_card_hbm_p5_arlock   ) ,
    .m_axi_card_hbm_p5_arprot       (m_axi_card_hbm_p5_arprot   ) ,
    .m_axi_card_hbm_p5_arqos        (m_axi_card_hbm_p5_arqos    ) ,
    .m_axi_card_hbm_p5_arready      (m_axi_card_hbm_p5_arready  ) ,
    .m_axi_card_hbm_p5_arregion     (m_axi_card_hbm_p5_arregion ) ,
    .m_axi_card_hbm_p5_arsize       (m_axi_card_hbm_p5_arsize   ) ,
    .m_axi_card_hbm_p5_aruser       (m_axi_card_hbm_p5_aruser   ) ,
    .m_axi_card_hbm_p5_arvalid      (m_axi_card_hbm_p5_arvalid  ) ,
    .m_axi_card_hbm_p5_awaddr       (temp_card_hbm_p5_awaddr    ) ,
    .m_axi_card_hbm_p5_awburst      (m_axi_card_hbm_p5_awburst  ) ,
    .m_axi_card_hbm_p5_awcache      (m_axi_card_hbm_p5_awcache  ) ,
    .m_axi_card_hbm_p5_awid         (m_axi_card_hbm_p5_awid     ) ,
    .m_axi_card_hbm_p5_awlen        (m_axi_card_hbm_p5_awlen    ) ,
    .m_axi_card_hbm_p5_awlock       (m_axi_card_hbm_p5_awlock   ) ,
    .m_axi_card_hbm_p5_awprot       (m_axi_card_hbm_p5_awprot   ) ,
    .m_axi_card_hbm_p5_awqos        (m_axi_card_hbm_p5_awqos    ) ,
    .m_axi_card_hbm_p5_awready      (m_axi_card_hbm_p5_awready  ) ,
    .m_axi_card_hbm_p5_awregion     (m_axi_card_hbm_p5_awregion ) ,
    .m_axi_card_hbm_p5_awsize       (m_axi_card_hbm_p5_awsize   ) ,
    .m_axi_card_hbm_p5_awuser       (m_axi_card_hbm_pp5awuser   ) ,
    .m_axi_card_hbm_p5_awvalid      (m_axi_card_hbm_p5_awvalid  ) ,
    .m_axi_card_hbm_p5_bid          (m_axi_card_hbm_p5_bid      ) ,
    .m_axi_card_hbm_p5_bready       (m_axi_card_hbm_p5_bready   ) ,
    .m_axi_card_hbm_p5_bresp        (m_axi_card_hbm_p5_bresp    ) ,
    .m_axi_card_hbm_p5_buser        (m_axi_card_hbm_p5_buser    ) ,
    .m_axi_card_hbm_p5_bvalid       (m_axi_card_hbm_p5_bvalid   ) ,
    .m_axi_card_hbm_p5_rdata        (m_axi_card_hbm_p5_rdata    ) ,
    .m_axi_card_hbm_p5_rid          (m_axi_card_hbm_p5_rid      ) ,
    .m_axi_card_hbm_p5_rlast        (m_axi_card_hbm_p5_rlast    ) ,
    .m_axi_card_hbm_p5_rready       (m_axi_card_hbm_p5_rready   ) ,
    .m_axi_card_hbm_p5_rresp        (m_axi_card_hbm_p5_rresp    ) ,
    .m_axi_card_hbm_p5_ruser        (m_axi_card_hbm_p5_ruser    ) ,
    .m_axi_card_hbm_p5_rvalid       (m_axi_card_hbm_p5_rvalid   ) ,
    .m_axi_card_hbm_p5_wdata        (m_axi_card_hbm_p5_wdata    ) ,
    .m_axi_card_hbm_p5_wid          (                           ) ,
    .m_axi_card_hbm_p5_wlast        (m_axi_card_hbm_p5_wlast    ) ,
    .m_axi_card_hbm_p5_wready       (m_axi_card_hbm_p5_wready   ) ,
    .m_axi_card_hbm_p5_wstrb        (m_axi_card_hbm_p5_wstrb    ) ,
    .m_axi_card_hbm_p5_wuser        (m_axi_card_hbm_p5_wuser    ) ,
    .m_axi_card_hbm_p5_wvalid       (m_axi_card_hbm_p5_wvalid   ) ,

    .m_axi_card_hbm_p6_araddr       (temp_card_hbm_p6_araddr    ) ,
    .m_axi_card_hbm_p6_arburst      (m_axi_card_hbm_p6_arburst  ) ,
    .m_axi_card_hbm_p6_arcache      (m_axi_card_hbm_p6_arcache  ) ,
    .m_axi_card_hbm_p6_arid         (m_axi_card_hbm_p6_arid     ) ,
    .m_axi_card_hbm_p6_arlen        (m_axi_card_hbm_p6_arlen    ) ,
    .m_axi_card_hbm_p6_arlock       (m_axi_card_hbm_p6_arlock   ) ,
    .m_axi_card_hbm_p6_arprot       (m_axi_card_hbm_p6_arprot   ) ,
    .m_axi_card_hbm_p6_arqos        (m_axi_card_hbm_p6_arqos    ) ,
    .m_axi_card_hbm_p6_arready      (m_axi_card_hbm_p6_arready  ) ,
    .m_axi_card_hbm_p6_arregion     (m_axi_card_hbm_p6_arregion ) ,
    .m_axi_card_hbm_p6_arsize       (m_axi_card_hbm_p6_arsize   ) ,
    .m_axi_card_hbm_p6_aruser       (m_axi_card_hbm_p6_aruser   ) ,
    .m_axi_card_hbm_p6_arvalid      (m_axi_card_hbm_p6_arvalid  ) ,
    .m_axi_card_hbm_p6_awaddr       (temp_card_hbm_p6_awaddr    ) ,
    .m_axi_card_hbm_p6_awburst      (m_axi_card_hbm_p6_awburst  ) ,
    .m_axi_card_hbm_p6_awcache      (m_axi_card_hbm_p6_awcache  ) ,
    .m_axi_card_hbm_p6_awid         (m_axi_card_hbm_p6_awid     ) ,
    .m_axi_card_hbm_p6_awlen        (m_axi_card_hbm_p6_awlen    ) ,
    .m_axi_card_hbm_p6_awlock       (m_axi_card_hbm_p6_awlock   ) ,
    .m_axi_card_hbm_p6_awprot       (m_axi_card_hbm_p6_awprot   ) ,
    .m_axi_card_hbm_p6_awqos        (m_axi_card_hbm_p6_awqos    ) ,
    .m_axi_card_hbm_p6_awready      (m_axi_card_hbm_p6_awready  ) ,
    .m_axi_card_hbm_p6_awregion     (m_axi_card_hbm_p6_awregion ) ,
    .m_axi_card_hbm_p6_awsize       (m_axi_card_hbm_p6_awsize   ) ,
    .m_axi_card_hbm_p6_awuser       (m_axi_card_hbm_p6_awuser   ) ,
    .m_axi_card_hbm_p6_awvalid      (m_axi_card_hbm_p6_awvalid  ) ,
    .m_axi_card_hbm_p6_bid          (m_axi_card_hbm_p6_bid      ) ,
    .m_axi_card_hbm_p6_bready       (m_axi_card_hbm_p6_bready   ) ,
    .m_axi_card_hbm_p6_bresp        (m_axi_card_hbm_p6_bresp    ) ,
    .m_axi_card_hbm_p6_buser        (m_axi_card_hbm_p6_buser    ) ,
    .m_axi_card_hbm_p6_bvalid       (m_axi_card_hbm_p6_bvalid   ) ,
    .m_axi_card_hbm_p6_rdata        (m_axi_card_hbm_p6_rdata    ) ,
    .m_axi_card_hbm_p6_rid          (m_axi_card_hbm_p6_rid      ) ,
    .m_axi_card_hbm_p6_rlast        (m_axi_card_hbm_p6_rlast    ) ,
    .m_axi_card_hbm_p6_rready       (m_axi_card_hbm_p6_rready   ) ,
    .m_axi_card_hbm_p6_rresp        (m_axi_card_hbm_p6_rresp    ) ,
    .m_axi_card_hbm_p6_ruser        (m_axi_card_hbm_p6_ruser    ) ,
    .m_axi_card_hbm_p6_rvalid       (m_axi_card_hbm_p6_rvalid   ) ,
    .m_axi_card_hbm_p6_wdata        (m_axi_card_hbm_p6_wdata    ) ,
    .m_axi_card_hbm_p6_wid          (                           ) ,
    .m_axi_card_hbm_p6_wlast        (m_axi_card_hbm_p6_wlast    ) ,
    .m_axi_card_hbm_p6_wready       (m_axi_card_hbm_p6_wready   ) ,
    .m_axi_card_hbm_p6_wstrb        (m_axi_card_hbm_p6_wstrb    ) ,
    .m_axi_card_hbm_p6_wuser        (m_axi_card_hbm_p6_wuser    ) ,
    .m_axi_card_hbm_p6_wvalid       (m_axi_card_hbm_p6_wvalid   ) ,

    .m_axi_card_hbm_p7_araddr       (temp_card_hbm_p7_araddr    ) ,
    .m_axi_card_hbm_p7_arburst      (m_axi_card_hbm_p7_arburst  ) ,
    .m_axi_card_hbm_p7_arcache      (m_axi_card_hbm_p7_arcache  ) ,
    .m_axi_card_hbm_p7_arid         (m_axi_card_hbm_p7_arid     ) ,
    .m_axi_card_hbm_p7_arlen        (m_axi_card_hbm_p7_arlen    ) ,
    .m_axi_card_hbm_p7_arlock       (m_axi_card_hbm_p7_arlock   ) ,
    .m_axi_card_hbm_p7_arprot       (m_axi_card_hbm_p7_arprot   ) ,
    .m_axi_card_hbm_p7_arqos        (m_axi_card_hbm_p7_arqos    ) ,
    .m_axi_card_hbm_p7_arready      (m_axi_card_hbm_p7_arready  ) ,
    .m_axi_card_hbm_p7_arregion     (m_axi_card_hbm_p7_arregion ) ,
    .m_axi_card_hbm_p7_arsize       (m_axi_card_hbm_p7_arsize   ) ,
    .m_axi_card_hbm_p7_aruser       (m_axi_card_hbm_p7_aruser   ) ,
    .m_axi_card_hbm_p7_arvalid      (m_axi_card_hbm_p7_arvalid  ) ,
    .m_axi_card_hbm_p7_awaddr       (temp_card_hbm_p7_awaddr    ) ,
    .m_axi_card_hbm_p7_awburst      (m_axi_card_hbm_p7_awburst  ) ,
    .m_axi_card_hbm_p7_awcache      (m_axi_card_hbm_p7_awcache  ) ,
    .m_axi_card_hbm_p7_awid         (m_axi_card_hbm_p7_awid     ) ,
    .m_axi_card_hbm_p7_awlen        (m_axi_card_hbm_p7_awlen    ) ,
    .m_axi_card_hbm_p7_awlock       (m_axi_card_hbm_p7_awlock   ) ,
    .m_axi_card_hbm_p7_awprot       (m_axi_card_hbm_p7_awprot   ) ,
    .m_axi_card_hbm_p7_awqos        (m_axi_card_hbm_p7_awqos    ) ,
    .m_axi_card_hbm_p7_awready      (m_axi_card_hbm_p7_awready  ) ,
    .m_axi_card_hbm_p7_awregion     (m_axi_card_hbm_p7_awregion ) ,
    .m_axi_card_hbm_p7_awsize       (m_axi_card_hbm_p7_awsize   ) ,
    .m_axi_card_hbm_p7_awuser       (m_axi_card_hbm_p7_awuser   ) ,
    .m_axi_card_hbm_p7_awvalid      (m_axi_card_hbm_p7_awvalid  ) ,
    .m_axi_card_hbm_p7_bid          (m_axi_card_hbm_p7_bid      ) ,
    .m_axi_card_hbm_p7_bready       (m_axi_card_hbm_p7_bready   ) ,
    .m_axi_card_hbm_p7_bresp        (m_axi_card_hbm_p7_bresp    ) ,
    .m_axi_card_hbm_p7_buser        (m_axi_card_hbm_p7_buser    ) ,
    .m_axi_card_hbm_p7_bvalid       (m_axi_card_hbm_p7_bvalid   ) ,
    .m_axi_card_hbm_p7_rdata        (m_axi_card_hbm_p7_rdata    ) ,
    .m_axi_card_hbm_p7_rid          (m_axi_card_hbm_p7_rid      ) ,
    .m_axi_card_hbm_p7_rlast        (m_axi_card_hbm_p7_rlast    ) ,
    .m_axi_card_hbm_p7_rready       (m_axi_card_hbm_p7_rready   ) ,
    .m_axi_card_hbm_p7_rresp        (m_axi_card_hbm_p7_rresp    ) ,
    .m_axi_card_hbm_p7_ruser        (m_axi_card_hbm_p7_ruser    ) ,
    .m_axi_card_hbm_p7_rvalid       (m_axi_card_hbm_p7_rvalid   ) ,
    .m_axi_card_hbm_p7_wdata        (m_axi_card_hbm_p7_wdata    ) ,
    .m_axi_card_hbm_p7_wid          (                           ) ,
    .m_axi_card_hbm_p7_wlast        (m_axi_card_hbm_p7_wlast    ) ,
    .m_axi_card_hbm_p7_wready       (m_axi_card_hbm_p7_wready   ) ,
    .m_axi_card_hbm_p7_wstrb        (m_axi_card_hbm_p7_wstrb    ) ,
    .m_axi_card_hbm_p7_wuser        (m_axi_card_hbm_p7_wuser    ) ,
    .m_axi_card_hbm_p7_wvalid       (m_axi_card_hbm_p7_wvalid   ) ,

    .m_axi_card_hbm_p8_araddr       (temp_card_hbm_p8_araddr    ) ,
    .m_axi_card_hbm_p8_arburst      (m_axi_card_hbm_p8_arburst  ) ,
    .m_axi_card_hbm_p8_arcache      (m_axi_card_hbm_p8_arcache  ) ,
    .m_axi_card_hbm_p8_arid         (m_axi_card_hbm_p8_arid     ) ,
    .m_axi_card_hbm_p8_arlen        (m_axi_card_hbm_p8_arlen    ) ,
    .m_axi_card_hbm_p8_arlock       (m_axi_card_hbm_p8_arlock   ) ,
    .m_axi_card_hbm_p8_arprot       (m_axi_card_hbm_p8_arprot   ) ,
    .m_axi_card_hbm_p8_arqos        (m_axi_card_hbm_p8_arqos    ) ,
    .m_axi_card_hbm_p8_arready      (m_axi_card_hbm_p8_arready  ) ,
    .m_axi_card_hbm_p8_arregion     (m_axi_card_hbm_p8_arregion ) ,
    .m_axi_card_hbm_p8_arsize       (m_axi_card_hbm_p8_arsize   ) ,
    .m_axi_card_hbm_p8_aruser       (m_axi_card_hbm_p8_aruser   ) ,
    .m_axi_card_hbm_p8_arvalid      (m_axi_card_hbm_p8_arvalid  ) ,
    .m_axi_card_hbm_p8_awaddr       (temp_card_hbm_p8_awaddr    ) ,
    .m_axi_card_hbm_p8_awburst      (m_axi_card_hbm_p8_awburst  ) ,
    .m_axi_card_hbm_p8_awcache      (m_axi_card_hbm_p8_awcache  ) ,
    .m_axi_card_hbm_p8_awid         (m_axi_card_hbm_p8_awid     ) ,
    .m_axi_card_hbm_p8_awlen        (m_axi_card_hbm_p8_awlen    ) ,
    .m_axi_card_hbm_p8_awlock       (m_axi_card_hbm_p8_awlock   ) ,
    .m_axi_card_hbm_p8_awprot       (m_axi_card_hbm_p8_awprot   ) ,
    .m_axi_card_hbm_p8_awqos        (m_axi_card_hbm_p8_awqos    ) ,
    .m_axi_card_hbm_p8_awready      (m_axi_card_hbm_p8_awready  ) ,
    .m_axi_card_hbm_p8_awregion     (m_axi_card_hbm_p8_awregion ) ,
    .m_axi_card_hbm_p8_awsize       (m_axi_card_hbm_p8_awsize   ) ,
    .m_axi_card_hbm_p8_awuser       (m_axi_card_hbm_p8_awuser   ) ,
    .m_axi_card_hbm_p8_awvalid      (m_axi_card_hbm_p8_awvalid  ) ,
    .m_axi_card_hbm_p8_bid          (m_axi_card_hbm_p8_bid      ) ,
    .m_axi_card_hbm_p8_bready       (m_axi_card_hbm_p8_bready   ) ,
    .m_axi_card_hbm_p8_bresp        (m_axi_card_hbm_p8_bresp    ) ,
    .m_axi_card_hbm_p8_buser        (m_axi_card_hbm_p8_buser    ) ,
    .m_axi_card_hbm_p8_bvalid       (m_axi_card_hbm_p8_bvalid   ) ,
    .m_axi_card_hbm_p8_rdata        (m_axi_card_hbm_p8_rdata    ) ,
    .m_axi_card_hbm_p8_rid          (m_axi_card_hbm_p8_rid      ) ,
    .m_axi_card_hbm_p8_rlast        (m_axi_card_hbm_p8_rlast    ) ,
    .m_axi_card_hbm_p8_rready       (m_axi_card_hbm_p8_rready   ) ,
    .m_axi_card_hbm_p8_rresp        (m_axi_card_hbm_p8_rresp    ) ,
    .m_axi_card_hbm_p8_ruser        (m_axi_card_hbm_p8_ruser    ) ,
    .m_axi_card_hbm_p8_rvalid       (m_axi_card_hbm_p8_rvalid   ) ,
    .m_axi_card_hbm_p8_wdata        (m_axi_card_hbm_p8_wdata    ) ,
    .m_axi_card_hbm_p8_wid          (                           ) ,
    .m_axi_card_hbm_p8_wlast        (m_axi_card_hbm_p8_wlast    ) ,
    .m_axi_card_hbm_p8_wready       (m_axi_card_hbm_p8_wready   ) ,
    .m_axi_card_hbm_p8_wstrb        (m_axi_card_hbm_p8_wstrb    ) ,
    .m_axi_card_hbm_p8_wuser        (m_axi_card_hbm_p8_wuser    ) ,
    .m_axi_card_hbm_p8_wvalid       (m_axi_card_hbm_p8_wvalid   ) ,

    .m_axi_card_hbm_p9_araddr       (temp_card_hbm_p9_araddr    ) ,
    .m_axi_card_hbm_p9_arburst      (m_axi_card_hbm_p9_arburst  ) ,
    .m_axi_card_hbm_p9_arcache      (m_axi_card_hbm_p9_arcache  ) ,
    .m_axi_card_hbm_p9_arid         (m_axi_card_hbm_p9_arid     ) ,
    .m_axi_card_hbm_p9_arlen        (m_axi_card_hbm_p9_arlen    ) ,
    .m_axi_card_hbm_p9_arlock       (m_axi_card_hbm_p9_arlock   ) ,
    .m_axi_card_hbm_p9_arprot       (m_axi_card_hbm_p9_arprot   ) ,
    .m_axi_card_hbm_p9_arqos        (m_axi_card_hbm_p9_arqos    ) ,
    .m_axi_card_hbm_p9_arready      (m_axi_card_hbm_p9_arready  ) ,
    .m_axi_card_hbm_p9_arregion     (m_axi_card_hbm_p9_arregion ) ,
    .m_axi_card_hbm_p9_arsize       (m_axi_card_hbm_p9_arsize   ) ,
    .m_axi_card_hbm_p9_aruser       (m_axi_card_hbm_p9_aruser   ) ,
    .m_axi_card_hbm_p9_arvalid      (m_axi_card_hbm_p9_arvalid  ) ,
    .m_axi_card_hbm_p9_awaddr       (temp_card_hbm_p9_awaddr    ) ,
    .m_axi_card_hbm_p9_awburst      (m_axi_card_hbm_p9_awburst  ) ,
    .m_axi_card_hbm_p9_awcache      (m_axi_card_hbm_p9_awcache  ) ,
    .m_axi_card_hbm_p9_awid         (m_axi_card_hbm_p9_awid     ) ,
    .m_axi_card_hbm_p9_awlen        (m_axi_card_hbm_p9_awlen    ) ,
    .m_axi_card_hbm_p9_awlock       (m_axi_card_hbm_p9_awlock   ) ,
    .m_axi_card_hbm_p9_awprot       (m_axi_card_hbm_p9_awprot   ) ,
    .m_axi_card_hbm_p9_awqos        (m_axi_card_hbm_p9_awqos    ) ,
    .m_axi_card_hbm_p9_awready      (m_axi_card_hbm_p9_awready  ) ,
    .m_axi_card_hbm_p9_awregion     (m_axi_card_hbm_p9_awregion ) ,
    .m_axi_card_hbm_p9_awsize       (m_axi_card_hbm_p9_awsize   ) ,
    .m_axi_card_hbm_p9_awuser       (m_axi_card_hbm_p9_awuser   ) ,
    .m_axi_card_hbm_p9_awvalid      (m_axi_card_hbm_p9_awvalid  ) ,
    .m_axi_card_hbm_p9_bid          (m_axi_card_hbm_p9_bid      ) ,
    .m_axi_card_hbm_p9_bready       (m_axi_card_hbm_p9_bready   ) ,
    .m_axi_card_hbm_p9_bresp        (m_axi_card_hbm_p9_bresp    ) ,
    .m_axi_card_hbm_p9_buser        (m_axi_card_hbm_p9_buser    ) ,
    .m_axi_card_hbm_p9_bvalid       (m_axi_card_hbm_p9_bvalid   ) ,
    .m_axi_card_hbm_p9_rdata        (m_axi_card_hbm_p9_rdata    ) ,
    .m_axi_card_hbm_p9_rid          (m_axi_card_hbm_p9_rid      ) ,
    .m_axi_card_hbm_p9_rlast        (m_axi_card_hbm_p9_rlast    ) ,
    .m_axi_card_hbm_p9_rready       (m_axi_card_hbm_p9_rready   ) ,
    .m_axi_card_hbm_p9_rresp        (m_axi_card_hbm_p9_rresp    ) ,
    .m_axi_card_hbm_p9_ruser        (m_axi_card_hbm_p9_ruser    ) ,
    .m_axi_card_hbm_p9_rvalid       (m_axi_card_hbm_p9_rvalid   ) ,
    .m_axi_card_hbm_p9_wdata        (m_axi_card_hbm_p9_wdata    ) ,
    .m_axi_card_hbm_p9_wid          (                           ) ,
    .m_axi_card_hbm_p9_wlast        (m_axi_card_hbm_p9_wlast    ) ,
    .m_axi_card_hbm_p9_wready       (m_axi_card_hbm_p9_wready   ) ,
    .m_axi_card_hbm_p9_wstrb        (m_axi_card_hbm_p9_wstrb    ) ,
    .m_axi_card_hbm_p9_wuser        (m_axi_card_hbm_p9_wuser    ) ,
    .m_axi_card_hbm_p9_wvalid       (m_axi_card_hbm_p9_wvalid   ) ,

    .m_axi_card_hbm_p10_araddr       (temp_card_hbm_p10_araddr    ) ,
    .m_axi_card_hbm_p10_arburst      (m_axi_card_hbm_p10_arburst  ) ,
    .m_axi_card_hbm_p10_arcache      (m_axi_card_hbm_p10_arcache  ) ,
    .m_axi_card_hbm_p10_arid         (m_axi_card_hbm_p10_arid     ) ,
    .m_axi_card_hbm_p10_arlen        (m_axi_card_hbm_p10_arlen    ) ,
    .m_axi_card_hbm_p10_arlock       (m_axi_card_hbm_p10_arlock   ) ,
    .m_axi_card_hbm_p10_arprot       (m_axi_card_hbm_p10_arprot   ) ,
    .m_axi_card_hbm_p10_arqos        (m_axi_card_hbm_p10_arqos    ) ,
    .m_axi_card_hbm_p10_arready      (m_axi_card_hbm_p10_arready  ) ,
    .m_axi_card_hbm_p10_arregion     (m_axi_card_hbm_p10_arregion ) ,
    .m_axi_card_hbm_p10_arsize       (m_axi_card_hbm_p10_arsize   ) ,
    .m_axi_card_hbm_p10_aruser       (m_axi_card_hbm_p10_aruser   ) ,
    .m_axi_card_hbm_p10_arvalid      (m_axi_card_hbm_p10_arvalid  ) ,
    .m_axi_card_hbm_p10_awaddr       (temp_card_hbm_p10_awaddr    ) ,
    .m_axi_card_hbm_p10_awburst      (m_axi_card_hbm_p10_awburst  ) ,
    .m_axi_card_hbm_p10_awcache      (m_axi_card_hbm_p10_awcache  ) ,
    .m_axi_card_hbm_p10_awid         (m_axi_card_hbm_p10_awid     ) ,
    .m_axi_card_hbm_p10_awlen        (m_axi_card_hbm_p10_awlen    ) ,
    .m_axi_card_hbm_p10_awlock       (m_axi_card_hbm_p10_awlock   ) ,
    .m_axi_card_hbm_p10_awprot       (m_axi_card_hbm_p10_awprot   ) ,
    .m_axi_card_hbm_p10_awqos        (m_axi_card_hbm_p10_awqos    ) ,
    .m_axi_card_hbm_p10_awready      (m_axi_card_hbm_p10_awready  ) ,
    .m_axi_card_hbm_p10_awregion     (m_axi_card_hbm_p10_awregion ) ,
    .m_axi_card_hbm_p10_awsize       (m_axi_card_hbm_p10_awsize   ) ,
    .m_axi_card_hbm_p10_awuser       (m_axi_card_hbm_p10_awuser   ) ,
    .m_axi_card_hbm_p10_awvalid      (m_axi_card_hbm_p10_awvalid  ) ,
    .m_axi_card_hbm_p10_bid          (m_axi_card_hbm_p10_bid      ) ,
    .m_axi_card_hbm_p10_bready       (m_axi_card_hbm_p10_bready   ) ,
    .m_axi_card_hbm_p10_bresp        (m_axi_card_hbm_p10_bresp    ) ,
    .m_axi_card_hbm_p10_buser        (m_axi_card_hbm_p10_buser    ) ,
    .m_axi_card_hbm_p10_bvalid       (m_axi_card_hbm_p10_bvalid   ) ,
    .m_axi_card_hbm_p10_rdata        (m_axi_card_hbm_p10_rdata    ) ,
    .m_axi_card_hbm_p10_rid          (m_axi_card_hbm_p10_rid      ) ,
    .m_axi_card_hbm_p10_rlast        (m_axi_card_hbm_p10_rlast    ) ,
    .m_axi_card_hbm_p10_rready       (m_axi_card_hbm_p10_rready   ) ,
    .m_axi_card_hbm_p10_rresp        (m_axi_card_hbm_p10_rresp    ) ,
    .m_axi_card_hbm_p10_ruser        (m_axi_card_hbm_p10_ruser    ) ,
    .m_axi_card_hbm_p10_rvalid       (m_axi_card_hbm_p10_rvalid   ) ,
    .m_axi_card_hbm_p10_wdata        (m_axi_card_hbm_p10_wdata    ) ,
    .m_axi_card_hbm_p10_wid          (                           ) ,
    .m_axi_card_hbm_p10_wlast        (m_axi_card_hbm_p10_wlast    ) ,
    .m_axi_card_hbm_p10_wready       (m_axi_card_hbm_p10_wready   ) ,
    .m_axi_card_hbm_p10_wstrb        (m_axi_card_hbm_p10_wstrb    ) ,
    .m_axi_card_hbm_p10_wuser        (m_axi_card_hbm_p10_wuser    ) ,
    .m_axi_card_hbm_p10_wvalid       (m_axi_card_hbm_p10_wvalid   ) ,

    .m_axi_card_hbm_p11_araddr       (temp_card_hbm_p11_araddr    ) ,
    .m_axi_card_hbm_p11_arburst      (m_axi_card_hbm_p11_arburst  ) ,
    .m_axi_card_hbm_p11_arcache      (m_axi_card_hbm_p11_arcache  ) ,
    .m_axi_card_hbm_p11_arid         (m_axi_card_hbm_p11_arid     ) ,
    .m_axi_card_hbm_p11_arlen        (m_axi_card_hbm_p11_arlen    ) ,
    .m_axi_card_hbm_p11_arlock       (m_axi_card_hbm_p11_arlock   ) ,
    .m_axi_card_hbm_p11_arprot       (m_axi_card_hbm_p11_arprot   ) ,
    .m_axi_card_hbm_p11_arqos        (m_axi_card_hbm_p11_arqos    ) ,
    .m_axi_card_hbm_p11_arready      (m_axi_card_hbm_p11_arready  ) ,
    .m_axi_card_hbm_p11_arregion     (m_axi_card_hbm_p11_arregion ) ,
    .m_axi_card_hbm_p11_arsize       (m_axi_card_hbm_p11_arsize   ) ,
    .m_axi_card_hbm_p11_aruser       (m_axi_card_hbm_p11_aruser   ) ,
    .m_axi_card_hbm_p11_arvalid      (m_axi_card_hbm_p11_arvalid  ) ,
    .m_axi_card_hbm_p11_awaddr       (temp_card_hbm_p11_awaddr    ) ,
    .m_axi_card_hbm_p11_awburst      (m_axi_card_hbm_p11_awburst  ) ,
    .m_axi_card_hbm_p11_awcache      (m_axi_card_hbm_p11_awcache  ) ,
    .m_axi_card_hbm_p11_awid         (m_axi_card_hbm_p11_awid     ) ,
    .m_axi_card_hbm_p11_awlen        (m_axi_card_hbm_p11_awlen    ) ,
    .m_axi_card_hbm_p11_awlock       (m_axi_card_hbm_p11_awlock   ) ,
    .m_axi_card_hbm_p11_awprot       (m_axi_card_hbm_p11_awprot   ) ,
    .m_axi_card_hbm_p11_awqos        (m_axi_card_hbm_p11_awqos    ) ,
    .m_axi_card_hbm_p11_awready      (m_axi_card_hbm_p11_awready  ) ,
    .m_axi_card_hbm_p11_awregion     (m_axi_card_hbm_p11_awregion ) ,
    .m_axi_card_hbm_p11_awsize       (m_axi_card_hbm_p11_awsize   ) ,
    .m_axi_card_hbm_p11_awuser       (m_axi_card_hbm_p11_awuser   ) ,
    .m_axi_card_hbm_p11_awvalid      (m_axi_card_hbm_p11_awvalid  ) ,
    .m_axi_card_hbm_p11_bid          (m_axi_card_hbm_p11_bid      ) ,
    .m_axi_card_hbm_p11_bready       (m_axi_card_hbm_p11_bready   ) ,
    .m_axi_card_hbm_p11_bresp        (m_axi_card_hbm_p11_bresp    ) ,
    .m_axi_card_hbm_p11_buser        (m_axi_card_hbm_p11_buser    ) ,
    .m_axi_card_hbm_p11_bvalid       (m_axi_card_hbm_p11_bvalid   ) ,
    .m_axi_card_hbm_p11_rdata        (m_axi_card_hbm_p11_rdata    ) ,
    .m_axi_card_hbm_p11_rid          (m_axi_card_hbm_p11_rid      ) ,
    .m_axi_card_hbm_p11_rlast        (m_axi_card_hbm_p11_rlast    ) ,
    .m_axi_card_hbm_p11_rready       (m_axi_card_hbm_p11_rready   ) ,
    .m_axi_card_hbm_p11_rresp        (m_axi_card_hbm_p11_rresp    ) ,
    .m_axi_card_hbm_p11_ruser        (m_axi_card_hbm_p11_ruser    ) ,
    .m_axi_card_hbm_p11_rvalid       (m_axi_card_hbm_p11_rvalid   ) ,
    .m_axi_card_hbm_p11_wdata        (m_axi_card_hbm_p11_wdata    ) ,
    .m_axi_card_hbm_p11_wid          (                           ) ,
    .m_axi_card_hbm_p11_wlast        (m_axi_card_hbm_p11_wlast    ) ,
    .m_axi_card_hbm_p11_wready       (m_axi_card_hbm_p11_wready   ) ,
    .m_axi_card_hbm_p11_wstrb        (m_axi_card_hbm_p11_wstrb    ) ,
    .m_axi_card_hbm_p11_wuser        (m_axi_card_hbm_p11_wuser    ) ,
    .m_axi_card_hbm_p11_wvalid       (m_axi_card_hbm_p11_wvalid   ) ,

`endif
`endif
    // ETHERNET interface
`ifdef ENABLE_ETHERNET
`ifndef ENABLE_ETH_LOOP_BACK
//ethernet enabled without loopback
    .din_eth_TDATA                (din_eth_TDATA            ) ,
    .din_eth_TVALID               (din_eth_TVALID           ) ,
    .din_eth_TREADY               (din_eth_TREADY           ) ,
    .din_eth_TKEEP                (din_eth_TKEEP            ) ,
    .din_eth_TUSER                (din_eth_TUSER            ) ,
    .din_eth_TLAST                (din_eth_TLAST            ) ,
//Enable for ethernet TX
    .dout_eth_TDATA               (dout_eth_TDATA           ) ,
    .dout_eth_TVALID              (dout_eth_TVALID          ) ,
    .dout_eth_TREADY              (dout_eth_TREADY          ) ,
    .dout_eth_TKEEP               (dout_eth_TKEEP           ) ,
    .dout_eth_TUSER               (dout_eth_TUSER           ) ,
    .dout_eth_TLAST               (dout_eth_TLAST           ) ,
    .eth_reset_V                  (eth_reset                ) ,
`else
    .din_eth_TDATA                (dwrap_eth_TDATA          ) ,
    .din_eth_TVALID               (dwrap_eth_TVALID         ) ,
    .din_eth_TREADY               (                         ) ,
    .din_eth_TKEEP                (dwrap_eth_TKEEP          ) ,
    .din_eth_TUSER                (dwrap_eth_TUSER          ) ,
    .din_eth_TLAST                (dwrap_eth_TLAST[0]       ) ,
//Enable for ethernet TX
    .dout_eth_TDATA               (dwrap_eth_TDATA          ) ,
    .dout_eth_TVALID              (dwrap_eth_TVALID         ) ,
//Force the TREADY signal to 1 to mimic the mac
    .dout_eth_TREADY              ('b1                      ) ,
    .dout_eth_TKEEP               (dwrap_eth_TKEEP          ) ,
    .dout_eth_TUSER               (dwrap_eth_TUSER          ) ,
    .dout_eth_TLAST               (dwrap_eth_TLAST[0]       ) ,
    .eth_reset_V                  (                         ) ,
//Enable ethernet with loopback
`endif
`endif
    //
    .s_axi_ctrl_reg_araddr        (s_axi_ctrl_reg_araddr    ) ,
    .s_axi_ctrl_reg_arready       (s_axi_ctrl_reg_arready   ) ,
    .s_axi_ctrl_reg_arvalid       (s_axi_ctrl_reg_arvalid   ) ,
    .s_axi_ctrl_reg_awaddr        (s_axi_ctrl_reg_awaddr    ) ,
    .s_axi_ctrl_reg_awready       (s_axi_ctrl_reg_awready   ) ,
    .s_axi_ctrl_reg_awvalid       (s_axi_ctrl_reg_awvalid   ) ,
    .s_axi_ctrl_reg_bready        (s_axi_ctrl_reg_bready    ) ,
    .s_axi_ctrl_reg_bresp         (s_axi_ctrl_reg_bresp     ) ,
    .s_axi_ctrl_reg_bvalid        (s_axi_ctrl_reg_bvalid    ) ,
    .s_axi_ctrl_reg_rdata         (temp_s_axi_ctrl_reg_rdata     ) ,
    .s_axi_ctrl_reg_rready        (s_axi_ctrl_reg_rready    ) ,
    .s_axi_ctrl_reg_rresp         (s_axi_ctrl_reg_rresp     ) ,
    .s_axi_ctrl_reg_rvalid        (s_axi_ctrl_reg_rvalid    ) ,
    .s_axi_ctrl_reg_wdata         (s_axi_ctrl_reg_wdata     ) ,
    .s_axi_ctrl_reg_wready        (s_axi_ctrl_reg_wready    ) ,
    .s_axi_ctrl_reg_wstrb         (s_axi_ctrl_reg_wstrb     ) ,
    .s_axi_ctrl_reg_wvalid        (s_axi_ctrl_reg_wvalid    ) ,
    .m_axi_host_mem_araddr        (m_axi_host_mem_araddr    ) ,
    .m_axi_host_mem_arburst       (m_axi_host_mem_arburst   ) ,
    .m_axi_host_mem_arcache       (m_axi_host_mem_arcache   ) ,
    .m_axi_host_mem_arid          (m_axi_host_mem_arid [0]  ) ,//SR# 10394170
    .m_axi_host_mem_arlen         (m_axi_host_mem_arlen     ) ,
    .m_axi_host_mem_arlock        (m_axi_host_mem_arlock    ) ,
    .m_axi_host_mem_arprot        (m_axi_host_mem_arprot    ) ,
    .m_axi_host_mem_arqos         (m_axi_host_mem_arqos     ) ,
    .m_axi_host_mem_arready       (m_axi_host_mem_arready   ) ,
    .m_axi_host_mem_arregion      (m_axi_host_mem_arregion  ) ,
    .m_axi_host_mem_arsize        (m_axi_host_mem_arsize    ) ,
    .m_axi_host_mem_aruser        (                         ) ,
    .m_axi_host_mem_arvalid       (m_axi_host_mem_arvalid   ) ,
    .m_axi_host_mem_awaddr        (m_axi_host_mem_awaddr    ) ,
    .m_axi_host_mem_awburst       (m_axi_host_mem_awburst   ) ,
    .m_axi_host_mem_awcache       (m_axi_host_mem_awcache   ) ,
    .m_axi_host_mem_awid          (m_axi_host_mem_awid [0]  ) ,//SR# 10394170
    .m_axi_host_mem_awlen         (m_axi_host_mem_awlen     ) ,
    .m_axi_host_mem_awlock        (m_axi_host_mem_awlock    ) ,
    .m_axi_host_mem_awprot        (m_axi_host_mem_awprot    ) ,
    .m_axi_host_mem_awqos         (m_axi_host_mem_awqos     ) ,
    .m_axi_host_mem_awready       (m_axi_host_mem_awready   ) ,
    .m_axi_host_mem_awregion      (m_axi_host_mem_awregion  ) ,
    .m_axi_host_mem_awsize        (m_axi_host_mem_awsize    ) ,
    .m_axi_host_mem_awuser        (                         ) ,
    .m_axi_host_mem_awvalid       (m_axi_host_mem_awvalid   ) ,
    .m_axi_host_mem_bid           (m_axi_host_mem_bid [0]   ) ,//SR# 10394170
    .m_axi_host_mem_bready        (m_axi_host_mem_bready    ) ,
    .m_axi_host_mem_bresp         (m_axi_host_mem_bresp     ) ,
    .m_axi_host_mem_buser         (m_axi_host_mem_buser [0] ) ,//SR# 10394170
    .m_axi_host_mem_bvalid        (m_axi_host_mem_bvalid    ) ,
    .m_axi_host_mem_rdata         (m_axi_host_mem_rdata     ) ,
    .m_axi_host_mem_rid           (m_axi_host_mem_rid [0]   ) ,//SR# 10394170
    .m_axi_host_mem_rlast         (m_axi_host_mem_rlast     ) ,
    .m_axi_host_mem_rready        (m_axi_host_mem_rready    ) ,
    .m_axi_host_mem_rresp         (m_axi_host_mem_rresp     ) ,
    .m_axi_host_mem_ruser         (m_axi_host_mem_ruser [0] ) ,//SR# 10394170
    .m_axi_host_mem_rvalid        (m_axi_host_mem_rvalid    ) ,
    .m_axi_host_mem_wdata         (m_axi_host_mem_wdata     ) ,
    .m_axi_host_mem_wid           (                         ) ,
    .m_axi_host_mem_wlast         (m_axi_host_mem_wlast     ) ,
    .m_axi_host_mem_wready        (m_axi_host_mem_wready    ) ,
    .m_axi_host_mem_wstrb         (m_axi_host_mem_wstrb     ) ,
    .m_axi_host_mem_wuser         (m_axi_host_mem_wuser [0] ) ,//SR# 10394170
    .m_axi_host_mem_wvalid        (m_axi_host_mem_wvalid    ) ,
    .interrupt                    ( interrupt_i             )
  );
//==========================================
// Reset for hls_action
always @ (posedge ap_clk)
     hls_rst_n_q <= ap_rst_n;

//==========================================
// Context is not implemented
always @ (posedge ap_clk)
    if (~ap_rst_n)
        context_q <= 0;
//    else if (s_axi_ctrl_reg_wvalid && (s_axi_ctrl_reg_awaddr = ADDR_CTX_ID_REG )
//        context_q <= s_axi_ctrl_reg_wdata;


//==========================================
// Interrupt handshaking logic
always @ (posedge ap_clk)
     if (~ap_rst_n) begin
        interrupt_q          <= 1'b0;
        interrupt_wait_ack_q <= 1'b0;
     end
     else begin
         interrupt_wait_ack_q <= (interrupt_i & ~interrupt_q ) | (interrupt_wait_ack_q & ~interrupt_ack);
         interrupt_q          <= interrupt_i & (interrupt_q | ~interrupt_wait_ack_q);
     end

// Interrupt output signals
  // Generating interrupt pulse
assign  interrupt     = interrupt_i & ~interrupt_q;
  // use fixed interrupt source id '0x4' for HLS interrupts
  // (the high order bit of the source id is assigned by SNAP)
always @ (posedge ap_clk)
    if (~ap_rst_n) begin
        interrupt_src_hi <= 32'b0;
        interrupt_src_lo <= 32'b0;
    end
    else if (s_axi_ctrl_reg_wvalid  && (s_axi_ctrl_reg_awaddr == ADDR_ACTION_INTERRUPT_SRC_ADDR_HI))
        interrupt_src_hi <= s_axi_ctrl_reg_wdata;
    else if (s_axi_ctrl_reg_wvalid  && (s_axi_ctrl_reg_awaddr == ADDR_ACTION_INTERRUPT_SRC_ADDR_LO))
        interrupt_src_lo <= s_axi_ctrl_reg_wdata;

assign  interrupt_src = {interrupt_src_hi, interrupt_src_lo};
  // context ID
assign  interrupt_ctx = context_q;


//==========================================
//When read ACTION_TYPE and RELEASE_LEVEL, the return data is handled here. 
//hls_action will return RVALID (acknowledgement), RDATA=0
//and RDATA is ORed with this reg_rdata_hijack. 
always @ (posedge ap_clk)
    if (~ap_rst_n) begin
        reg_rdata_hijack <= 32'h0;
    end
    else if (s_axi_ctrl_reg_arvalid == 1'b1) begin
        if (s_axi_ctrl_reg_araddr == ADDR_ACTION_TYPE)
            reg_rdata_hijack <= `HLS_ACTION_TYPE;
        else if (s_axi_ctrl_reg_araddr == ADDR_RELEASE_LEVEL)
            reg_rdata_hijack <= `HLS_RELEASE_LEVEL;
        else
            reg_rdata_hijack <= 32'h0;
    end

assign s_axi_ctrl_reg_rdata = reg_rdata_hijack | temp_s_axi_ctrl_reg_rdata;

//==========================================
// Driving context ID to host memory interface
assign  m_axi_host_mem_aruser = context_q;
assign  m_axi_host_mem_awuser = context_q;

// Driving the higher ID fields to 0.
generate if(`IDW > 1)
begin:high_hid_fields_driver
    assign  m_axi_host_mem_arid  [ `IDW-1 : 1 ] = 'b0;
    assign  m_axi_host_mem_awid  [ `IDW-1 : 1 ] = 'b0;
end
endgenerate
//assign  m_axi_host_mem_wuser [ `AXI_WUSER-1 : 1 ] = 'b0;


// if DDR or DDR replaced by BRAM
`ifdef ENABLE_AXI_CARD_MEM
`ifndef ENABLE_HBM
assign m_axi_card_mem0_araddr = temp_card_mem0_araddr[`AXI_CARD_MEM_ADDR_WIDTH-1:0];
assign m_axi_card_mem0_awaddr = temp_card_mem0_awaddr[`AXI_CARD_MEM_ADDR_WIDTH-1:0];

generate if(`AXI_CARD_MEM_ID_WIDTH > 1)
begin:high_cid_fields_driver
    assign m_axi_card_mem0_arid  [ `AXI_CARD_MEM_ID_WIDTH-1 : 1 ] = 'b0;
    assign m_axi_card_mem0_awid  [ `AXI_CARD_MEM_ID_WIDTH-1 : 1 ] = 'b0;
end
endgenerate

// if HBM
`else
assign m_axi_card_hbm_p0_araddr = temp_card_hbm_p0_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p0_awaddr = temp_card_hbm_p0_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p1_araddr = temp_card_hbm_p1_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p1_awaddr = temp_card_hbm_p1_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p2_araddr = temp_card_hbm_p2_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p2_awaddr = temp_card_hbm_p2_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p3_araddr = temp_card_hbm_p3_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p3_awaddr = temp_card_hbm_p3_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p4_araddr = temp_card_hbm_p4_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p4_awaddr = temp_card_hbm_p4_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p5_araddr = temp_card_hbm_p5_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p5_awaddr = temp_card_hbm_p5_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p6_araddr = temp_card_hbm_p6_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p6_awaddr = temp_card_hbm_p6_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p7_araddr = temp_card_hbm_p7_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p7_awaddr = temp_card_hbm_p7_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p8_araddr = temp_card_hbm_p8_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p8_awaddr = temp_card_hbm_p8_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p9_araddr = temp_card_hbm_p9_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p9_awaddr = temp_card_hbm_p9_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p10_araddr = temp_card_hbm_p10_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p10_awaddr = temp_card_hbm_p10_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p11_araddr = temp_card_hbm_p11_araddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];
assign m_axi_card_hbm_p11_awaddr = temp_card_hbm_p11_awaddr[`AXI_CARD_HBM_ADDR_WIDTH-1:0];

`endif
`endif
endmodule
