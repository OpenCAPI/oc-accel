// *********************************************************************
// IBM CONFIDENTIAL BACKGROUND TECHNOLOGY: VERIFICATION ENVIRONMENT FILE
// *********************************************************************

`ifndef _SB_SVH
`define _SB_SVH


`include "tl_mem_model.sv"
`include "tl_scoreboard.sv"

`endif

