`ifndef _TL_BFM_PKG_SVH_
`define _TL_BFM_PKG_SVH_

//CONFIG
//INTERFACE & TRANSACTIONS
//MANAGER
`include "../util/util.svh"

//SCOREBOARDS
`include "../sb/sb.svh"

//MONITORS
//DRIVER
//AGENTS
`include "../tl/tl.svh"

//TL BFM TOP
//`include "tl_bfm_env.sv"

//TEST LIST
`include "../seq_lib/test_list.svh"

`endif // _TL_BFM_PKG_SVH_
