// *********************************************************************
// IBM CONFIDENTIAL BACKGROUND TECHNOLOGY: VERIFICATION ENVIRONMENT FILE
// *********************************************************************

`ifndef _TEST_LIST_SVH
`define _TEST_LIST_SVH

`include "bfm_sequence_base.sv"
`include "bfm_seq_lib.sv"
`include "bfm_seq_lib_rand_resp.sv"
`include "bfm_seq_lib_rand_axi.sv"
`include "bfm_seq_lib_rand_axi_resp.sv"
`include "odma_seq_lib.sv"
`include "odma_seq_lib_unalign.sv"
`include "bfm_seq_lib_mmio_intrp.sv"

`endif
